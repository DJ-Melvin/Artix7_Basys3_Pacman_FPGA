`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////
// Module Name: get_font
/////////////////////////////////////////////////////////////////

// font.coe
module get_font(
    input [13:0] addr,
    output reg [11:0] color
);  
    always@(*) begin
        case(addr)
            0: color = 12'h000;
            1: color = 12'h000;
            2: color = 12'h000;
            3: color = 12'h000;
            4: color = 12'h000;
            5: color = 12'h000;
            6: color = 12'h000;
            7: color = 12'h000;
            8: color = 12'h000;
            9: color = 12'h000;
            10: color = 12'h000;
            11: color = 12'h000;
            12: color = 12'h000;
            13: color = 12'h000;
            14: color = 12'h000;
            15: color = 12'h000;
            16: color = 12'h000;
            17: color = 12'h000;
            18: color = 12'h000;
            19: color = 12'h000;
            20: color = 12'h000;
            21: color = 12'h000;
            22: color = 12'h000;
            23: color = 12'h000;
            24: color = 12'h000;
            25: color = 12'h000;
            26: color = 12'h000;
            27: color = 12'h000;
            28: color = 12'h000;
            29: color = 12'h000;
            30: color = 12'h000;
            31: color = 12'h000;
            32: color = 12'h000;
            33: color = 12'h000;
            34: color = 12'h000;
            35: color = 12'h000;
            36: color = 12'h000;
            37: color = 12'h000;
            38: color = 12'h000;
            39: color = 12'h000;
            40: color = 12'h000;
            41: color = 12'h000;
            42: color = 12'h000;
            43: color = 12'h000;
            44: color = 12'h000;
            45: color = 12'h000;
            46: color = 12'h000;
            47: color = 12'h000;
            48: color = 12'h000;
            49: color = 12'h000;
            50: color = 12'h000;
            51: color = 12'h000;
            52: color = 12'h000;
            53: color = 12'h000;
            54: color = 12'h000;
            55: color = 12'h000;
            56: color = 12'h000;
            57: color = 12'h000;
            58: color = 12'h000;
            59: color = 12'h000;
            60: color = 12'h000;
            61: color = 12'h000;
            62: color = 12'h000;
            63: color = 12'h000;
            64: color = 12'h000;
            65: color = 12'h000;
            66: color = 12'h000;
            67: color = 12'h000;
            68: color = 12'h000;
            69: color = 12'h000;
            70: color = 12'h000;
            71: color = 12'h000;
            72: color = 12'h000;
            73: color = 12'h000;
            74: color = 12'h000;
            75: color = 12'h000;
            76: color = 12'h000;
            77: color = 12'h000;
            78: color = 12'h000;
            79: color = 12'h000;
            80: color = 12'h000;
            81: color = 12'h000;
            82: color = 12'h000;
            83: color = 12'h000;
            84: color = 12'h000;
            85: color = 12'h000;
            86: color = 12'h000;
            87: color = 12'h000;
            88: color = 12'h000;
            89: color = 12'h000;
            90: color = 12'h000;
            91: color = 12'h000;
            92: color = 12'h000;
            93: color = 12'h000;
            94: color = 12'h000;
            95: color = 12'h000;
            96: color = 12'h000;
            97: color = 12'h000;
            98: color = 12'h000;
            99: color = 12'h000;
            100: color = 12'h000;
            101: color = 12'h000;
            102: color = 12'h000;
            103: color = 12'h000;
            104: color = 12'h000;
            105: color = 12'h000;
            106: color = 12'h000;
            107: color = 12'h000;
            108: color = 12'h000;
            109: color = 12'h000;
            110: color = 12'h000;
            111: color = 12'h000;
            112: color = 12'h000;
            113: color = 12'h000;
            114: color = 12'h000;
            115: color = 12'h000;
            116: color = 12'h000;
            117: color = 12'h000;
            118: color = 12'h000;
            119: color = 12'h000;
            120: color = 12'h000;
            121: color = 12'h000;
            122: color = 12'h000;
            123: color = 12'h000;
            124: color = 12'h000;
            125: color = 12'h000;
            126: color = 12'h000;
            127: color = 12'h000;
            128: color = 12'h000;
            129: color = 12'h000;
            130: color = 12'h000;
            131: color = 12'h000;
            132: color = 12'h000;
            133: color = 12'h000;
            134: color = 12'h000;
            135: color = 12'h000;
            136: color = 12'h000;
            137: color = 12'h000;
            138: color = 12'h000;
            139: color = 12'h000;
            140: color = 12'h000;
            141: color = 12'h000;
            142: color = 12'h000;
            143: color = 12'h000;
            144: color = 12'h000;
            145: color = 12'h000;
            146: color = 12'h000;
            147: color = 12'h000;
            148: color = 12'h000;
            149: color = 12'h000;
            150: color = 12'h000;
            151: color = 12'h000;
            152: color = 12'h000;
            153: color = 12'h000;
            154: color = 12'h000;
            155: color = 12'h000;
            156: color = 12'h000;
            157: color = 12'h000;
            158: color = 12'h000;
            159: color = 12'h000;
            160: color = 12'h000;
            161: color = 12'h000;
            162: color = 12'h000;
            163: color = 12'h000;
            164: color = 12'h000;
            165: color = 12'h000;
            166: color = 12'h000;
            167: color = 12'h000;
            168: color = 12'h000;
            169: color = 12'h000;
            170: color = 12'h000;
            171: color = 12'h000;
            172: color = 12'h000;
            173: color = 12'h000;
            174: color = 12'h000;
            175: color = 12'h000;
            176: color = 12'h000;
            177: color = 12'h000;
            178: color = 12'h000;
            179: color = 12'h000;
            180: color = 12'h000;
            181: color = 12'h000;
            182: color = 12'h000;
            183: color = 12'h000;
            184: color = 12'h000;
            185: color = 12'h000;
            186: color = 12'h000;
            187: color = 12'h000;
            188: color = 12'h000;
            189: color = 12'h000;
            190: color = 12'h000;
            191: color = 12'h000;
            192: color = 12'h000;
            193: color = 12'h000;
            194: color = 12'h000;
            195: color = 12'h000;
            196: color = 12'h000;
            197: color = 12'h000;
            198: color = 12'h000;
            199: color = 12'h000;
            200: color = 12'h000;
            201: color = 12'h000;
            202: color = 12'h000;
            203: color = 12'h000;
            204: color = 12'h000;
            205: color = 12'h000;
            206: color = 12'h000;
            207: color = 12'h000;
            208: color = 12'h000;
            209: color = 12'h000;
            210: color = 12'h000;
            211: color = 12'h000;
            212: color = 12'h000;
            213: color = 12'h000;
            214: color = 12'h000;
            215: color = 12'h000;
            216: color = 12'h000;
            217: color = 12'h000;
            218: color = 12'h000;
            219: color = 12'h000;
            220: color = 12'h000;
            221: color = 12'h000;
            222: color = 12'h000;
            223: color = 12'h000;
            224: color = 12'h000;
            225: color = 12'h000;
            226: color = 12'h000;
            227: color = 12'h000;
            228: color = 12'h000;
            229: color = 12'h000;
            230: color = 12'h000;
            231: color = 12'h000;
            232: color = 12'h000;
            233: color = 12'h000;
            234: color = 12'h000;
            235: color = 12'h000;
            236: color = 12'h000;
            237: color = 12'h000;
            238: color = 12'h000;
            239: color = 12'h000;
            240: color = 12'h000;
            241: color = 12'h000;
            242: color = 12'h000;
            243: color = 12'h000;
            244: color = 12'h000;
            245: color = 12'h000;
            246: color = 12'h000;
            247: color = 12'h000;
            248: color = 12'h000;
            249: color = 12'h000;
            250: color = 12'h000;
            251: color = 12'h000;
            252: color = 12'h000;
            253: color = 12'h000;
            254: color = 12'h000;
            255: color = 12'h000;
            256: color = 12'h000;
            257: color = 12'h000;
            258: color = 12'h000;
            259: color = 12'h000;
            260: color = 12'h000;
            261: color = 12'h000;
            262: color = 12'h000;
            263: color = 12'h000;
            264: color = 12'h000;
            265: color = 12'h000;
            266: color = 12'h000;
            267: color = 12'h000;
            268: color = 12'h000;
            269: color = 12'h000;
            270: color = 12'h000;
            271: color = 12'h000;
            272: color = 12'h000;
            273: color = 12'h000;
            274: color = 12'h000;
            275: color = 12'h000;
            276: color = 12'h000;
            277: color = 12'h000;
            278: color = 12'h000;
            279: color = 12'h000;
            280: color = 12'h000;
            281: color = 12'h000;
            282: color = 12'h000;
            283: color = 12'h000;
            284: color = 12'h000;
            285: color = 12'h000;
            286: color = 12'h000;
            287: color = 12'h000;
            288: color = 12'h000;
            289: color = 12'h000;
            290: color = 12'h000;
            291: color = 12'h000;
            292: color = 12'h000;
            293: color = 12'h000;
            294: color = 12'h000;
            295: color = 12'h000;
            296: color = 12'h000;
            297: color = 12'h000;
            298: color = 12'h000;
            299: color = 12'h000;
            300: color = 12'h000;
            301: color = 12'h000;
            302: color = 12'h000;
            303: color = 12'h000;
            304: color = 12'h000;
            305: color = 12'h000;
            306: color = 12'h000;
            307: color = 12'h000;
            308: color = 12'h000;
            309: color = 12'h000;
            310: color = 12'h000;
            311: color = 12'h000;
            312: color = 12'h000;
            313: color = 12'h000;
            314: color = 12'h000;
            315: color = 12'h000;
            316: color = 12'h000;
            317: color = 12'h000;
            318: color = 12'h000;
            319: color = 12'h000;
            320: color = 12'h000;
            321: color = 12'h000;
            322: color = 12'h000;
            323: color = 12'h000;
            324: color = 12'h000;
            325: color = 12'h000;
            326: color = 12'h000;
            327: color = 12'h000;
            328: color = 12'h000;
            329: color = 12'h000;
            330: color = 12'h000;
            331: color = 12'h000;
            332: color = 12'h000;
            333: color = 12'h000;
            334: color = 12'h000;
            335: color = 12'h000;
            336: color = 12'h000;
            337: color = 12'h000;
            338: color = 12'h000;
            339: color = 12'h000;
            340: color = 12'h000;
            341: color = 12'h000;
            342: color = 12'h000;
            343: color = 12'h000;
            344: color = 12'h000;
            345: color = 12'h000;
            346: color = 12'h000;
            347: color = 12'h000;
            348: color = 12'h000;
            349: color = 12'h000;
            350: color = 12'h000;
            351: color = 12'h000;
            352: color = 12'h000;
            353: color = 12'h000;
            354: color = 12'h000;
            355: color = 12'h000;
            356: color = 12'h000;
            357: color = 12'h000;
            358: color = 12'h000;
            359: color = 12'h000;
            360: color = 12'h000;
            361: color = 12'h000;
            362: color = 12'h000;
            363: color = 12'h000;
            364: color = 12'h000;
            365: color = 12'h000;
            366: color = 12'h000;
            367: color = 12'h000;
            368: color = 12'h000;
            369: color = 12'h000;
            370: color = 12'h000;
            371: color = 12'h000;
            372: color = 12'h000;
            373: color = 12'h000;
            374: color = 12'h000;
            375: color = 12'h000;
            376: color = 12'h000;
            377: color = 12'h000;
            378: color = 12'h000;
            379: color = 12'h000;
            380: color = 12'h000;
            381: color = 12'h000;
            382: color = 12'h000;
            383: color = 12'h000;
            384: color = 12'h000;
            385: color = 12'h000;
            386: color = 12'h000;
            387: color = 12'h000;
            388: color = 12'h000;
            389: color = 12'h000;
            390: color = 12'h000;
            391: color = 12'h000;
            392: color = 12'h000;
            393: color = 12'h000;
            394: color = 12'h000;
            395: color = 12'h000;
            396: color = 12'h000;
            397: color = 12'h000;
            398: color = 12'h000;
            399: color = 12'h000;
            400: color = 12'h000;
            401: color = 12'h000;
            402: color = 12'h000;
            403: color = 12'h000;
            404: color = 12'h000;
            405: color = 12'h000;
            406: color = 12'h000;
            407: color = 12'h000;
            408: color = 12'h000;
            409: color = 12'h000;
            410: color = 12'h000;
            411: color = 12'h000;
            412: color = 12'h000;
            413: color = 12'h000;
            414: color = 12'h000;
            415: color = 12'h000;
            416: color = 12'h000;
            417: color = 12'h000;
            418: color = 12'h000;
            419: color = 12'h000;
            420: color = 12'h000;
            421: color = 12'h000;
            422: color = 12'h000;
            423: color = 12'h000;
            424: color = 12'h000;
            425: color = 12'h000;
            426: color = 12'h000;
            427: color = 12'h000;
            428: color = 12'h000;
            429: color = 12'h000;
            430: color = 12'h000;
            431: color = 12'h000;
            432: color = 12'h000;
            433: color = 12'h000;
            434: color = 12'h000;
            435: color = 12'h000;
            436: color = 12'h000;
            437: color = 12'h000;
            438: color = 12'h000;
            439: color = 12'h000;
            440: color = 12'h000;
            441: color = 12'h000;
            442: color = 12'h000;
            443: color = 12'h000;
            444: color = 12'h000;
            445: color = 12'h000;
            446: color = 12'h000;
            447: color = 12'h000;
            448: color = 12'h000;
            449: color = 12'h000;
            450: color = 12'h000;
            451: color = 12'h000;
            452: color = 12'h000;
            453: color = 12'h000;
            454: color = 12'h000;
            455: color = 12'h000;
            456: color = 12'h000;
            457: color = 12'h000;
            458: color = 12'h000;
            459: color = 12'h000;
            460: color = 12'h000;
            461: color = 12'h000;
            462: color = 12'h000;
            463: color = 12'h000;
            464: color = 12'h000;
            465: color = 12'h000;
            466: color = 12'h000;
            467: color = 12'h000;
            468: color = 12'h000;
            469: color = 12'h000;
            470: color = 12'h000;
            471: color = 12'h000;
            472: color = 12'h000;
            473: color = 12'h000;
            474: color = 12'h000;
            475: color = 12'h000;
            476: color = 12'h000;
            477: color = 12'h000;
            478: color = 12'h000;
            479: color = 12'h000;
            480: color = 12'h000;
            481: color = 12'h000;
            482: color = 12'h000;
            483: color = 12'h000;
            484: color = 12'h000;
            485: color = 12'h000;
            486: color = 12'h000;
            487: color = 12'h000;
            488: color = 12'h000;
            489: color = 12'h000;
            490: color = 12'h000;
            491: color = 12'h000;
            492: color = 12'h000;
            493: color = 12'h000;
            494: color = 12'h000;
            495: color = 12'h000;
            496: color = 12'h000;
            497: color = 12'h000;
            498: color = 12'h000;
            499: color = 12'h000;
            500: color = 12'h000;
            501: color = 12'h000;
            502: color = 12'h000;
            503: color = 12'h000;
            504: color = 12'h000;
            505: color = 12'h000;
            506: color = 12'h000;
            507: color = 12'h000;
            508: color = 12'h000;
            509: color = 12'h000;
            510: color = 12'h000;
            511: color = 12'h000;
            512: color = 12'h000;
            513: color = 12'h000;
            514: color = 12'h000;
            515: color = 12'h000;
            516: color = 12'h000;
            517: color = 12'h000;
            518: color = 12'h000;
            519: color = 12'h000;
            520: color = 12'h000;
            521: color = 12'h000;
            522: color = 12'h000;
            523: color = 12'h000;
            524: color = 12'h000;
            525: color = 12'h000;
            526: color = 12'h000;
            527: color = 12'h000;
            528: color = 12'h000;
            529: color = 12'h000;
            530: color = 12'h000;
            531: color = 12'h000;
            532: color = 12'h000;
            533: color = 12'h000;
            534: color = 12'h000;
            535: color = 12'h000;
            536: color = 12'h000;
            537: color = 12'h000;
            538: color = 12'h000;
            539: color = 12'h000;
            540: color = 12'h000;
            541: color = 12'h000;
            542: color = 12'h000;
            543: color = 12'h000;
            544: color = 12'h000;
            545: color = 12'h000;
            546: color = 12'h000;
            547: color = 12'h000;
            548: color = 12'h000;
            549: color = 12'h000;
            550: color = 12'h000;
            551: color = 12'h000;
            552: color = 12'h000;
            553: color = 12'h000;
            554: color = 12'h000;
            555: color = 12'h000;
            556: color = 12'h000;
            557: color = 12'h000;
            558: color = 12'h000;
            559: color = 12'h000;
            560: color = 12'h000;
            561: color = 12'h000;
            562: color = 12'h000;
            563: color = 12'h000;
            564: color = 12'h000;
            565: color = 12'h000;
            566: color = 12'h000;
            567: color = 12'h000;
            568: color = 12'h000;
            569: color = 12'h000;
            570: color = 12'h000;
            571: color = 12'h000;
            572: color = 12'h000;
            573: color = 12'h000;
            574: color = 12'h000;
            575: color = 12'h000;
            576: color = 12'h000;
            577: color = 12'h000;
            578: color = 12'h000;
            579: color = 12'h000;
            580: color = 12'h000;
            581: color = 12'h000;
            582: color = 12'h000;
            583: color = 12'h000;
            584: color = 12'h000;
            585: color = 12'h000;
            586: color = 12'h000;
            587: color = 12'h000;
            588: color = 12'h000;
            589: color = 12'h000;
            590: color = 12'h000;
            591: color = 12'h000;
            592: color = 12'h000;
            593: color = 12'h000;
            594: color = 12'h000;
            595: color = 12'h000;
            596: color = 12'h000;
            597: color = 12'h000;
            598: color = 12'h000;
            599: color = 12'h000;
            600: color = 12'h000;
            601: color = 12'h000;
            602: color = 12'h000;
            603: color = 12'h000;
            604: color = 12'h000;
            605: color = 12'h000;
            606: color = 12'h000;
            607: color = 12'h000;
            608: color = 12'h000;
            609: color = 12'h000;
            610: color = 12'h000;
            611: color = 12'h000;
            612: color = 12'h000;
            613: color = 12'h000;
            614: color = 12'h000;
            615: color = 12'h000;
            616: color = 12'h000;
            617: color = 12'h000;
            618: color = 12'h000;
            619: color = 12'h000;
            620: color = 12'h000;
            621: color = 12'h000;
            622: color = 12'h000;
            623: color = 12'h000;
            624: color = 12'h000;
            625: color = 12'h000;
            626: color = 12'h000;
            627: color = 12'h000;
            628: color = 12'h000;
            629: color = 12'h000;
            630: color = 12'h000;
            631: color = 12'h000;
            632: color = 12'h000;
            633: color = 12'h000;
            634: color = 12'h000;
            635: color = 12'h000;
            636: color = 12'h000;
            637: color = 12'h000;
            638: color = 12'h000;
            639: color = 12'h000;
            640: color = 12'h000;
            641: color = 12'h000;
            642: color = 12'h000;
            643: color = 12'h000;
            644: color = 12'h000;
            645: color = 12'h000;
            646: color = 12'h000;
            647: color = 12'h000;
            648: color = 12'h000;
            649: color = 12'h000;
            650: color = 12'h000;
            651: color = 12'h000;
            652: color = 12'h000;
            653: color = 12'h000;
            654: color = 12'h000;
            655: color = 12'h000;
            656: color = 12'h000;
            657: color = 12'h000;
            658: color = 12'h000;
            659: color = 12'h000;
            660: color = 12'h000;
            661: color = 12'h000;
            662: color = 12'h000;
            663: color = 12'h000;
            664: color = 12'h000;
            665: color = 12'h000;
            666: color = 12'h000;
            667: color = 12'h000;
            668: color = 12'h000;
            669: color = 12'h000;
            670: color = 12'h000;
            671: color = 12'h000;
            672: color = 12'h000;
            673: color = 12'h000;
            674: color = 12'h000;
            675: color = 12'h000;
            676: color = 12'h000;
            677: color = 12'h000;
            678: color = 12'h000;
            679: color = 12'h000;
            680: color = 12'h000;
            681: color = 12'h000;
            682: color = 12'h000;
            683: color = 12'h000;
            684: color = 12'h000;
            685: color = 12'h000;
            686: color = 12'h000;
            687: color = 12'h000;
            688: color = 12'h000;
            689: color = 12'h000;
            690: color = 12'h000;
            691: color = 12'h000;
            692: color = 12'h000;
            693: color = 12'h000;
            694: color = 12'h000;
            695: color = 12'h000;
            696: color = 12'h000;
            697: color = 12'h000;
            698: color = 12'h000;
            699: color = 12'h000;
            700: color = 12'h000;
            701: color = 12'h000;
            702: color = 12'h000;
            703: color = 12'h000;
            704: color = 12'h000;
            705: color = 12'h000;
            706: color = 12'h000;
            707: color = 12'h000;
            708: color = 12'h000;
            709: color = 12'h000;
            710: color = 12'h000;
            711: color = 12'h000;
            712: color = 12'h000;
            713: color = 12'h000;
            714: color = 12'h000;
            715: color = 12'h000;
            716: color = 12'h000;
            717: color = 12'h000;
            718: color = 12'h000;
            719: color = 12'h000;
            720: color = 12'h000;
            721: color = 12'h000;
            722: color = 12'h000;
            723: color = 12'h000;
            724: color = 12'h000;
            725: color = 12'h000;
            726: color = 12'h000;
            727: color = 12'h000;
            728: color = 12'h000;
            729: color = 12'h000;
            730: color = 12'h000;
            731: color = 12'h000;
            732: color = 12'h000;
            733: color = 12'h000;
            734: color = 12'h000;
            735: color = 12'h000;
            736: color = 12'h000;
            737: color = 12'h000;
            738: color = 12'h000;
            739: color = 12'h000;
            740: color = 12'h000;
            741: color = 12'h000;
            742: color = 12'h000;
            743: color = 12'h000;
            744: color = 12'h000;
            745: color = 12'h000;
            746: color = 12'h000;
            747: color = 12'h000;
            748: color = 12'h000;
            749: color = 12'h000;
            750: color = 12'h000;
            751: color = 12'h000;
            752: color = 12'h000;
            753: color = 12'h000;
            754: color = 12'h000;
            755: color = 12'h000;
            756: color = 12'h000;
            757: color = 12'h000;
            758: color = 12'h000;
            759: color = 12'h000;
            760: color = 12'h000;
            761: color = 12'h000;
            762: color = 12'h000;
            763: color = 12'h000;
            764: color = 12'h000;
            765: color = 12'h000;
            766: color = 12'h000;
            767: color = 12'h000;
            768: color = 12'h000;
            769: color = 12'h000;
            770: color = 12'h000;
            771: color = 12'h000;
            772: color = 12'h000;
            773: color = 12'h000;
            774: color = 12'h000;
            775: color = 12'h000;
            776: color = 12'h000;
            777: color = 12'h000;
            778: color = 12'h000;
            779: color = 12'h000;
            780: color = 12'h000;
            781: color = 12'h000;
            782: color = 12'h000;
            783: color = 12'h000;
            784: color = 12'h000;
            785: color = 12'h000;
            786: color = 12'h000;
            787: color = 12'h000;
            788: color = 12'h000;
            789: color = 12'h000;
            790: color = 12'h000;
            791: color = 12'h000;
            792: color = 12'h000;
            793: color = 12'h000;
            794: color = 12'h000;
            795: color = 12'h000;
            796: color = 12'h000;
            797: color = 12'h000;
            798: color = 12'h000;
            799: color = 12'h000;
            800: color = 12'h000;
            801: color = 12'h000;
            802: color = 12'h000;
            803: color = 12'h000;
            804: color = 12'h000;
            805: color = 12'h000;
            806: color = 12'h000;
            807: color = 12'h000;
            808: color = 12'h000;
            809: color = 12'h000;
            810: color = 12'h000;
            811: color = 12'h000;
            812: color = 12'h000;
            813: color = 12'h000;
            814: color = 12'h000;
            815: color = 12'h000;
            816: color = 12'h000;
            817: color = 12'h000;
            818: color = 12'h000;
            819: color = 12'h000;
            820: color = 12'h000;
            821: color = 12'h000;
            822: color = 12'h000;
            823: color = 12'h000;
            824: color = 12'h000;
            825: color = 12'h000;
            826: color = 12'h000;
            827: color = 12'h000;
            828: color = 12'h000;
            829: color = 12'h000;
            830: color = 12'h000;
            831: color = 12'h000;
            832: color = 12'h000;
            833: color = 12'h000;
            834: color = 12'h000;
            835: color = 12'h000;
            836: color = 12'h000;
            837: color = 12'h000;
            838: color = 12'h000;
            839: color = 12'h000;
            840: color = 12'h000;
            841: color = 12'h000;
            842: color = 12'h000;
            843: color = 12'h000;
            844: color = 12'h000;
            845: color = 12'h000;
            846: color = 12'h000;
            847: color = 12'h000;
            848: color = 12'h000;
            849: color = 12'h000;
            850: color = 12'h000;
            851: color = 12'h000;
            852: color = 12'h000;
            853: color = 12'h000;
            854: color = 12'h000;
            855: color = 12'h000;
            856: color = 12'h000;
            857: color = 12'h000;
            858: color = 12'h000;
            859: color = 12'h000;
            860: color = 12'h000;
            861: color = 12'h000;
            862: color = 12'h000;
            863: color = 12'h000;
            864: color = 12'h000;
            865: color = 12'h000;
            866: color = 12'h000;
            867: color = 12'h000;
            868: color = 12'h000;
            869: color = 12'h000;
            870: color = 12'h000;
            871: color = 12'h000;
            872: color = 12'h000;
            873: color = 12'h000;
            874: color = 12'h000;
            875: color = 12'h000;
            876: color = 12'h000;
            877: color = 12'h000;
            878: color = 12'h000;
            879: color = 12'h000;
            880: color = 12'h000;
            881: color = 12'h000;
            882: color = 12'h000;
            883: color = 12'h000;
            884: color = 12'h000;
            885: color = 12'h000;
            886: color = 12'h000;
            887: color = 12'h000;
            888: color = 12'h000;
            889: color = 12'h000;
            890: color = 12'h000;
            891: color = 12'h000;
            892: color = 12'h000;
            893: color = 12'h000;
            894: color = 12'h000;
            895: color = 12'h000;
            896: color = 12'h000;
            897: color = 12'h000;
            898: color = 12'h000;
            899: color = 12'h000;
            900: color = 12'h000;
            901: color = 12'h000;
            902: color = 12'h000;
            903: color = 12'h000;
            904: color = 12'h000;
            905: color = 12'h000;
            906: color = 12'h000;
            907: color = 12'h000;
            908: color = 12'h000;
            909: color = 12'h000;
            910: color = 12'h000;
            911: color = 12'h000;
            912: color = 12'h000;
            913: color = 12'h000;
            914: color = 12'h000;
            915: color = 12'h000;
            916: color = 12'h000;
            917: color = 12'h000;
            918: color = 12'h000;
            919: color = 12'h000;
            920: color = 12'h000;
            921: color = 12'h000;
            922: color = 12'h000;
            923: color = 12'h000;
            924: color = 12'h000;
            925: color = 12'h000;
            926: color = 12'h000;
            927: color = 12'h000;
            928: color = 12'h000;
            929: color = 12'h000;
            930: color = 12'h000;
            931: color = 12'h000;
            932: color = 12'h000;
            933: color = 12'h000;
            934: color = 12'h000;
            935: color = 12'h000;
            936: color = 12'h000;
            937: color = 12'h000;
            938: color = 12'h000;
            939: color = 12'h000;
            940: color = 12'h000;
            941: color = 12'h000;
            942: color = 12'h000;
            943: color = 12'h000;
            944: color = 12'h000;
            945: color = 12'h000;
            946: color = 12'h000;
            947: color = 12'h000;
            948: color = 12'h000;
            949: color = 12'h000;
            950: color = 12'h000;
            951: color = 12'h000;
            952: color = 12'h000;
            953: color = 12'h000;
            954: color = 12'h000;
            955: color = 12'h000;
            956: color = 12'h000;
            957: color = 12'h000;
            958: color = 12'h000;
            959: color = 12'h000;
            960: color = 12'h000;
            961: color = 12'h000;
            962: color = 12'h000;
            963: color = 12'h000;
            964: color = 12'h000;
            965: color = 12'h000;
            966: color = 12'h000;
            967: color = 12'h000;
            968: color = 12'h000;
            969: color = 12'h000;
            970: color = 12'h000;
            971: color = 12'h000;
            972: color = 12'h000;
            973: color = 12'h000;
            974: color = 12'h000;
            975: color = 12'h000;
            976: color = 12'h000;
            977: color = 12'h000;
            978: color = 12'h000;
            979: color = 12'h000;
            980: color = 12'h000;
            981: color = 12'h000;
            982: color = 12'h000;
            983: color = 12'h000;
            984: color = 12'h000;
            985: color = 12'h000;
            986: color = 12'h000;
            987: color = 12'h000;
            988: color = 12'h000;
            989: color = 12'h000;
            990: color = 12'h000;
            991: color = 12'h000;
            992: color = 12'h000;
            993: color = 12'h000;
            994: color = 12'h000;
            995: color = 12'h000;
            996: color = 12'h000;
            997: color = 12'h000;
            998: color = 12'h000;
            999: color = 12'h000;
            1000: color = 12'h000;
            1001: color = 12'h000;
            1002: color = 12'h000;
            1003: color = 12'h000;
            1004: color = 12'h000;
            1005: color = 12'h000;
            1006: color = 12'h000;
            1007: color = 12'h000;
            1008: color = 12'h000;
            1009: color = 12'h000;
            1010: color = 12'h000;
            1011: color = 12'h000;
            1012: color = 12'h000;
            1013: color = 12'h000;
            1014: color = 12'h000;
            1015: color = 12'h000;
            1016: color = 12'h000;
            1017: color = 12'h000;
            1018: color = 12'h000;
            1019: color = 12'h000;
            1020: color = 12'h000;
            1021: color = 12'h000;
            1022: color = 12'h000;
            1023: color = 12'h000;
            1024: color = 12'h000;
            1025: color = 12'h000;
            1026: color = 12'h000;
            1027: color = 12'h000;
            1028: color = 12'h000;
            1029: color = 12'h000;
            1030: color = 12'h000;
            1031: color = 12'h000;
            1032: color = 12'h000;
            1033: color = 12'h000;
            1034: color = 12'h000;
            1035: color = 12'h000;
            1036: color = 12'h000;
            1037: color = 12'h000;
            1038: color = 12'h000;
            1039: color = 12'h000;
            1040: color = 12'h000;
            1041: color = 12'h000;
            1042: color = 12'h000;
            1043: color = 12'h000;
            1044: color = 12'h000;
            1045: color = 12'h000;
            1046: color = 12'h000;
            1047: color = 12'h000;
            1048: color = 12'h000;
            1049: color = 12'h000;
            1050: color = 12'h000;
            1051: color = 12'h000;
            1052: color = 12'h000;
            1053: color = 12'h000;
            1054: color = 12'h000;
            1055: color = 12'h000;
            1056: color = 12'h000;
            1057: color = 12'h000;
            1058: color = 12'h000;
            1059: color = 12'h000;
            1060: color = 12'h000;
            1061: color = 12'h000;
            1062: color = 12'h000;
            1063: color = 12'h000;
            1064: color = 12'h000;
            1065: color = 12'h000;
            1066: color = 12'h000;
            1067: color = 12'h000;
            1068: color = 12'h000;
            1069: color = 12'h000;
            1070: color = 12'h000;
            1071: color = 12'h000;
            1072: color = 12'h000;
            1073: color = 12'h000;
            1074: color = 12'h000;
            1075: color = 12'h000;
            1076: color = 12'h000;
            1077: color = 12'h000;
            1078: color = 12'h000;
            1079: color = 12'h000;
            1080: color = 12'h000;
            1081: color = 12'h000;
            1082: color = 12'h000;
            1083: color = 12'h000;
            1084: color = 12'h000;
            1085: color = 12'h000;
            1086: color = 12'h000;
            1087: color = 12'h000;
            1088: color = 12'h000;
            1089: color = 12'h000;
            1090: color = 12'h000;
            1091: color = 12'h000;
            1092: color = 12'h000;
            1093: color = 12'h000;
            1094: color = 12'h000;
            1095: color = 12'h000;
            1096: color = 12'h000;
            1097: color = 12'h000;
            1098: color = 12'h000;
            1099: color = 12'h000;
            1100: color = 12'h000;
            1101: color = 12'h000;
            1102: color = 12'h000;
            1103: color = 12'h000;
            1104: color = 12'h000;
            1105: color = 12'h000;
            1106: color = 12'h000;
            1107: color = 12'h000;
            1108: color = 12'h000;
            1109: color = 12'h000;
            1110: color = 12'h000;
            1111: color = 12'h000;
            1112: color = 12'h000;
            1113: color = 12'h000;
            1114: color = 12'h000;
            1115: color = 12'h000;
            1116: color = 12'h000;
            1117: color = 12'h000;
            1118: color = 12'h000;
            1119: color = 12'h000;
            1120: color = 12'h000;
            1121: color = 12'h000;
            1122: color = 12'h000;
            1123: color = 12'h000;
            1124: color = 12'h000;
            1125: color = 12'h000;
            1126: color = 12'h000;
            1127: color = 12'h000;
            1128: color = 12'h000;
            1129: color = 12'h000;
            1130: color = 12'h000;
            1131: color = 12'h000;
            1132: color = 12'h000;
            1133: color = 12'h000;
            1134: color = 12'h000;
            1135: color = 12'h000;
            1136: color = 12'h000;
            1137: color = 12'h000;
            1138: color = 12'h000;
            1139: color = 12'h000;
            1140: color = 12'h000;
            1141: color = 12'h000;
            1142: color = 12'h000;
            1143: color = 12'h000;
            1144: color = 12'h000;
            1145: color = 12'h000;
            1146: color = 12'h000;
            1147: color = 12'h000;
            1148: color = 12'h000;
            1149: color = 12'h000;
            1150: color = 12'h000;
            1151: color = 12'h000;
            1152: color = 12'h000;
            1153: color = 12'h000;
            1154: color = 12'h000;
            1155: color = 12'h000;
            1156: color = 12'h000;
            1157: color = 12'h000;
            1158: color = 12'h000;
            1159: color = 12'h000;
            1160: color = 12'h000;
            1161: color = 12'h000;
            1162: color = 12'h000;
            1163: color = 12'h000;
            1164: color = 12'h000;
            1165: color = 12'h000;
            1166: color = 12'h000;
            1167: color = 12'h000;
            1168: color = 12'h000;
            1169: color = 12'h000;
            1170: color = 12'h000;
            1171: color = 12'h000;
            1172: color = 12'h000;
            1173: color = 12'h000;
            1174: color = 12'h000;
            1175: color = 12'h000;
            1176: color = 12'h000;
            1177: color = 12'h000;
            1178: color = 12'h000;
            1179: color = 12'h000;
            1180: color = 12'h000;
            1181: color = 12'h000;
            1182: color = 12'h000;
            1183: color = 12'h000;
            1184: color = 12'h000;
            1185: color = 12'h000;
            1186: color = 12'h000;
            1187: color = 12'h000;
            1188: color = 12'h000;
            1189: color = 12'h000;
            1190: color = 12'h000;
            1191: color = 12'h000;
            1192: color = 12'h000;
            1193: color = 12'h000;
            1194: color = 12'h000;
            1195: color = 12'h000;
            1196: color = 12'h000;
            1197: color = 12'h000;
            1198: color = 12'h000;
            1199: color = 12'h000;
            1200: color = 12'h000;
            1201: color = 12'h000;
            1202: color = 12'h000;
            1203: color = 12'h000;
            1204: color = 12'h000;
            1205: color = 12'h000;
            1206: color = 12'h000;
            1207: color = 12'h000;
            1208: color = 12'h000;
            1209: color = 12'h000;
            1210: color = 12'h000;
            1211: color = 12'h000;
            1212: color = 12'h000;
            1213: color = 12'h000;
            1214: color = 12'h000;
            1215: color = 12'h000;
            1216: color = 12'h000;
            1217: color = 12'h000;
            1218: color = 12'h000;
            1219: color = 12'h000;
            1220: color = 12'h000;
            1221: color = 12'h000;
            1222: color = 12'h000;
            1223: color = 12'h000;
            1224: color = 12'h000;
            1225: color = 12'h000;
            1226: color = 12'h000;
            1227: color = 12'h000;
            1228: color = 12'h000;
            1229: color = 12'h000;
            1230: color = 12'h000;
            1231: color = 12'h000;
            1232: color = 12'h000;
            1233: color = 12'h000;
            1234: color = 12'h000;
            1235: color = 12'h000;
            1236: color = 12'h000;
            1237: color = 12'h000;
            1238: color = 12'h000;
            1239: color = 12'h000;
            1240: color = 12'h000;
            1241: color = 12'h000;
            1242: color = 12'h000;
            1243: color = 12'h000;
            1244: color = 12'h000;
            1245: color = 12'h000;
            1246: color = 12'h000;
            1247: color = 12'h000;
            1248: color = 12'h000;
            1249: color = 12'h000;
            1250: color = 12'h000;
            1251: color = 12'h000;
            1252: color = 12'h000;
            1253: color = 12'h000;
            1254: color = 12'h000;
            1255: color = 12'h000;
            1256: color = 12'h000;
            1257: color = 12'h000;
            1258: color = 12'h000;
            1259: color = 12'h000;
            1260: color = 12'h000;
            1261: color = 12'h000;
            1262: color = 12'h000;
            1263: color = 12'h000;
            1264: color = 12'h000;
            1265: color = 12'h000;
            1266: color = 12'h000;
            1267: color = 12'h000;
            1268: color = 12'h000;
            1269: color = 12'h000;
            1270: color = 12'h000;
            1271: color = 12'h000;
            1272: color = 12'h000;
            1273: color = 12'h000;
            1274: color = 12'h000;
            1275: color = 12'h000;
            1276: color = 12'h000;
            1277: color = 12'h000;
            1278: color = 12'h000;
            1279: color = 12'h000;
            1280: color = 12'h000;
            1281: color = 12'h000;
            1282: color = 12'h000;
            1283: color = 12'h000;
            1284: color = 12'h000;
            1285: color = 12'h000;
            1286: color = 12'h000;
            1287: color = 12'h000;
            1288: color = 12'h000;
            1289: color = 12'h000;
            1290: color = 12'h000;
            1291: color = 12'h000;
            1292: color = 12'h000;
            1293: color = 12'h000;
            1294: color = 12'h000;
            1295: color = 12'h000;
            1296: color = 12'h000;
            1297: color = 12'h000;
            1298: color = 12'h000;
            1299: color = 12'h000;
            1300: color = 12'h000;
            1301: color = 12'h000;
            1302: color = 12'h000;
            1303: color = 12'h000;
            1304: color = 12'h000;
            1305: color = 12'h000;
            1306: color = 12'h000;
            1307: color = 12'h000;
            1308: color = 12'h000;
            1309: color = 12'h000;
            1310: color = 12'h000;
            1311: color = 12'h000;
            1312: color = 12'h000;
            1313: color = 12'h000;
            1314: color = 12'h000;
            1315: color = 12'h000;
            1316: color = 12'h000;
            1317: color = 12'h000;
            1318: color = 12'h000;
            1319: color = 12'h000;
            1320: color = 12'h000;
            1321: color = 12'h000;
            1322: color = 12'h000;
            1323: color = 12'h000;
            1324: color = 12'h000;
            1325: color = 12'h000;
            1326: color = 12'h000;
            1327: color = 12'h000;
            1328: color = 12'h000;
            1329: color = 12'h000;
            1330: color = 12'h000;
            1331: color = 12'h000;
            1332: color = 12'h000;
            1333: color = 12'h000;
            1334: color = 12'h000;
            1335: color = 12'h000;
            1336: color = 12'h000;
            1337: color = 12'h000;
            1338: color = 12'h000;
            1339: color = 12'h000;
            1340: color = 12'h000;
            1341: color = 12'h000;
            1342: color = 12'h000;
            1343: color = 12'h000;
            1344: color = 12'h000;
            1345: color = 12'h000;
            1346: color = 12'h000;
            1347: color = 12'h000;
            1348: color = 12'h000;
            1349: color = 12'h000;
            1350: color = 12'h000;
            1351: color = 12'h000;
            1352: color = 12'h000;
            1353: color = 12'h000;
            1354: color = 12'h000;
            1355: color = 12'h000;
            1356: color = 12'h000;
            1357: color = 12'h000;
            1358: color = 12'h000;
            1359: color = 12'h000;
            1360: color = 12'h000;
            1361: color = 12'h000;
            1362: color = 12'h000;
            1363: color = 12'h000;
            1364: color = 12'h000;
            1365: color = 12'h000;
            1366: color = 12'h000;
            1367: color = 12'h000;
            1368: color = 12'h000;
            1369: color = 12'h000;
            1370: color = 12'h000;
            1371: color = 12'h000;
            1372: color = 12'h000;
            1373: color = 12'h000;
            1374: color = 12'h000;
            1375: color = 12'h000;
            1376: color = 12'h000;
            1377: color = 12'h000;
            1378: color = 12'h000;
            1379: color = 12'h000;
            1380: color = 12'h000;
            1381: color = 12'h000;
            1382: color = 12'h000;
            1383: color = 12'h000;
            1384: color = 12'h000;
            1385: color = 12'h000;
            1386: color = 12'h000;
            1387: color = 12'h000;
            1388: color = 12'h000;
            1389: color = 12'h000;
            1390: color = 12'h000;
            1391: color = 12'h000;
            1392: color = 12'h000;
            1393: color = 12'h000;
            1394: color = 12'h000;
            1395: color = 12'h000;
            1396: color = 12'h000;
            1397: color = 12'h000;
            1398: color = 12'h000;
            1399: color = 12'h000;
            1400: color = 12'h000;
            1401: color = 12'h000;
            1402: color = 12'h000;
            1403: color = 12'h000;
            1404: color = 12'h000;
            1405: color = 12'h000;
            1406: color = 12'h000;
            1407: color = 12'h000;
            1408: color = 12'h000;
            1409: color = 12'h000;
            1410: color = 12'h000;
            1411: color = 12'h000;
            1412: color = 12'h000;
            1413: color = 12'h000;
            1414: color = 12'h000;
            1415: color = 12'h000;
            1416: color = 12'h000;
            1417: color = 12'h000;
            1418: color = 12'h000;
            1419: color = 12'h000;
            1420: color = 12'h000;
            1421: color = 12'h000;
            1422: color = 12'h000;
            1423: color = 12'h000;
            1424: color = 12'h000;
            1425: color = 12'h000;
            1426: color = 12'h000;
            1427: color = 12'h000;
            1428: color = 12'h000;
            1429: color = 12'h000;
            1430: color = 12'h000;
            1431: color = 12'h000;
            1432: color = 12'h000;
            1433: color = 12'h000;
            1434: color = 12'h000;
            1435: color = 12'h000;
            1436: color = 12'h000;
            1437: color = 12'h000;
            1438: color = 12'h000;
            1439: color = 12'h000;
            1440: color = 12'h000;
            1441: color = 12'h000;
            1442: color = 12'h000;
            1443: color = 12'h000;
            1444: color = 12'h000;
            1445: color = 12'h000;
            1446: color = 12'h000;
            1447: color = 12'h000;
            1448: color = 12'h000;
            1449: color = 12'h000;
            1450: color = 12'h000;
            1451: color = 12'h000;
            1452: color = 12'h000;
            1453: color = 12'h000;
            1454: color = 12'h000;
            1455: color = 12'h000;
            1456: color = 12'h000;
            1457: color = 12'h000;
            1458: color = 12'h000;
            1459: color = 12'h000;
            1460: color = 12'h000;
            1461: color = 12'h000;
            1462: color = 12'h000;
            1463: color = 12'h000;
            1464: color = 12'h000;
            1465: color = 12'h000;
            1466: color = 12'h000;
            1467: color = 12'h000;
            1468: color = 12'h000;
            1469: color = 12'h000;
            1470: color = 12'h000;
            1471: color = 12'h000;
            1472: color = 12'h000;
            1473: color = 12'h000;
            1474: color = 12'h000;
            1475: color = 12'h000;
            1476: color = 12'h000;
            1477: color = 12'h000;
            1478: color = 12'h000;
            1479: color = 12'h000;
            1480: color = 12'h000;
            1481: color = 12'h000;
            1482: color = 12'h000;
            1483: color = 12'h000;
            1484: color = 12'h000;
            1485: color = 12'h000;
            1486: color = 12'h000;
            1487: color = 12'h000;
            1488: color = 12'h000;
            1489: color = 12'h000;
            1490: color = 12'h000;
            1491: color = 12'h000;
            1492: color = 12'h000;
            1493: color = 12'h000;
            1494: color = 12'h000;
            1495: color = 12'h000;
            1496: color = 12'h000;
            1497: color = 12'h000;
            1498: color = 12'h000;
            1499: color = 12'h000;
            1500: color = 12'h000;
            1501: color = 12'h000;
            1502: color = 12'h000;
            1503: color = 12'h000;
            1504: color = 12'h000;
            1505: color = 12'h000;
            1506: color = 12'h000;
            1507: color = 12'h000;
            1508: color = 12'h000;
            1509: color = 12'h000;
            1510: color = 12'h000;
            1511: color = 12'h000;
            1512: color = 12'h000;
            1513: color = 12'h000;
            1514: color = 12'h000;
            1515: color = 12'h000;
            1516: color = 12'h000;
            1517: color = 12'h000;
            1518: color = 12'h000;
            1519: color = 12'h000;
            1520: color = 12'h000;
            1521: color = 12'h000;
            1522: color = 12'h000;
            1523: color = 12'h000;
            1524: color = 12'h000;
            1525: color = 12'h000;
            1526: color = 12'h000;
            1527: color = 12'h000;
            1528: color = 12'h000;
            1529: color = 12'h000;
            1530: color = 12'h000;
            1531: color = 12'h000;
            1532: color = 12'h000;
            1533: color = 12'h000;
            1534: color = 12'h000;
            1535: color = 12'h000;
            1536: color = 12'h000;
            1537: color = 12'h000;
            1538: color = 12'h000;
            1539: color = 12'h000;
            1540: color = 12'h000;
            1541: color = 12'h000;
            1542: color = 12'h000;
            1543: color = 12'h000;
            1544: color = 12'h000;
            1545: color = 12'h000;
            1546: color = 12'h000;
            1547: color = 12'h000;
            1548: color = 12'h000;
            1549: color = 12'h000;
            1550: color = 12'h000;
            1551: color = 12'h000;
            1552: color = 12'h000;
            1553: color = 12'h000;
            1554: color = 12'h000;
            1555: color = 12'h000;
            1556: color = 12'h000;
            1557: color = 12'h000;
            1558: color = 12'h000;
            1559: color = 12'h000;
            1560: color = 12'h000;
            1561: color = 12'h000;
            1562: color = 12'h000;
            1563: color = 12'h000;
            1564: color = 12'h000;
            1565: color = 12'h000;
            1566: color = 12'h000;
            1567: color = 12'h000;
            1568: color = 12'h000;
            1569: color = 12'h000;
            1570: color = 12'h000;
            1571: color = 12'h000;
            1572: color = 12'h000;
            1573: color = 12'h000;
            1574: color = 12'h000;
            1575: color = 12'h000;
            1576: color = 12'h000;
            1577: color = 12'h000;
            1578: color = 12'h000;
            1579: color = 12'h000;
            1580: color = 12'h000;
            1581: color = 12'h000;
            1582: color = 12'h000;
            1583: color = 12'h000;
            1584: color = 12'h000;
            1585: color = 12'h000;
            1586: color = 12'h000;
            1587: color = 12'h000;
            1588: color = 12'h000;
            1589: color = 12'h000;
            1590: color = 12'h000;
            1591: color = 12'h000;
            1592: color = 12'h000;
            1593: color = 12'h000;
            1594: color = 12'h000;
            1595: color = 12'h000;
            1596: color = 12'h000;
            1597: color = 12'h000;
            1598: color = 12'h000;
            1599: color = 12'h000;
            1600: color = 12'h000;
            1601: color = 12'h000;
            1602: color = 12'h000;
            1603: color = 12'h000;
            1604: color = 12'h000;
            1605: color = 12'h000;
            1606: color = 12'h000;
            1607: color = 12'h000;
            1608: color = 12'h000;
            1609: color = 12'h000;
            1610: color = 12'h000;
            1611: color = 12'h000;
            1612: color = 12'h000;
            1613: color = 12'h000;
            1614: color = 12'h000;
            1615: color = 12'h000;
            1616: color = 12'h000;
            1617: color = 12'h000;
            1618: color = 12'h000;
            1619: color = 12'h000;
            1620: color = 12'h000;
            1621: color = 12'h000;
            1622: color = 12'h000;
            1623: color = 12'h000;
            1624: color = 12'h000;
            1625: color = 12'h000;
            1626: color = 12'h000;
            1627: color = 12'h000;
            1628: color = 12'h000;
            1629: color = 12'h000;
            1630: color = 12'h000;
            1631: color = 12'h000;
            1632: color = 12'h000;
            1633: color = 12'h000;
            1634: color = 12'h000;
            1635: color = 12'h000;
            1636: color = 12'h000;
            1637: color = 12'h000;
            1638: color = 12'h000;
            1639: color = 12'h000;
            1640: color = 12'h000;
            1641: color = 12'h000;
            1642: color = 12'h000;
            1643: color = 12'h000;
            1644: color = 12'h000;
            1645: color = 12'h000;
            1646: color = 12'h000;
            1647: color = 12'h000;
            1648: color = 12'h000;
            1649: color = 12'h000;
            1650: color = 12'h000;
            1651: color = 12'h000;
            1652: color = 12'h000;
            1653: color = 12'h000;
            1654: color = 12'h000;
            1655: color = 12'h000;
            1656: color = 12'h000;
            1657: color = 12'h000;
            1658: color = 12'h000;
            1659: color = 12'h000;
            1660: color = 12'h000;
            1661: color = 12'h000;
            1662: color = 12'h000;
            1663: color = 12'h000;
            1664: color = 12'h000;
            1665: color = 12'h000;
            1666: color = 12'h000;
            1667: color = 12'h000;
            1668: color = 12'h000;
            1669: color = 12'h000;
            1670: color = 12'h000;
            1671: color = 12'h000;
            1672: color = 12'h000;
            1673: color = 12'h000;
            1674: color = 12'h000;
            1675: color = 12'h000;
            1676: color = 12'h000;
            1677: color = 12'h000;
            1678: color = 12'h000;
            1679: color = 12'h000;
            1680: color = 12'h000;
            1681: color = 12'h000;
            1682: color = 12'h000;
            1683: color = 12'h000;
            1684: color = 12'h000;
            1685: color = 12'h000;
            1686: color = 12'h000;
            1687: color = 12'h000;
            1688: color = 12'h000;
            1689: color = 12'h000;
            1690: color = 12'h000;
            1691: color = 12'h000;
            1692: color = 12'h000;
            1693: color = 12'h000;
            1694: color = 12'h000;
            1695: color = 12'h000;
            1696: color = 12'h000;
            1697: color = 12'h000;
            1698: color = 12'h000;
            1699: color = 12'h000;
            1700: color = 12'h000;
            1701: color = 12'h000;
            1702: color = 12'h000;
            1703: color = 12'h000;
            1704: color = 12'h000;
            1705: color = 12'h000;
            1706: color = 12'h000;
            1707: color = 12'h000;
            1708: color = 12'h000;
            1709: color = 12'h000;
            1710: color = 12'h000;
            1711: color = 12'h000;
            1712: color = 12'h000;
            1713: color = 12'h000;
            1714: color = 12'h000;
            1715: color = 12'h000;
            1716: color = 12'h000;
            1717: color = 12'h000;
            1718: color = 12'h000;
            1719: color = 12'h000;
            1720: color = 12'h000;
            1721: color = 12'h000;
            1722: color = 12'h000;
            1723: color = 12'h000;
            1724: color = 12'h000;
            1725: color = 12'h000;
            1726: color = 12'h000;
            1727: color = 12'h000;
            1728: color = 12'h000;
            1729: color = 12'h000;
            1730: color = 12'h000;
            1731: color = 12'h000;
            1732: color = 12'h000;
            1733: color = 12'h000;
            1734: color = 12'h000;
            1735: color = 12'h000;
            1736: color = 12'h000;
            1737: color = 12'h000;
            1738: color = 12'h000;
            1739: color = 12'h000;
            1740: color = 12'h000;
            1741: color = 12'h000;
            1742: color = 12'h000;
            1743: color = 12'h000;
            1744: color = 12'h000;
            1745: color = 12'h000;
            1746: color = 12'h000;
            1747: color = 12'h000;
            1748: color = 12'h000;
            1749: color = 12'h000;
            1750: color = 12'h000;
            1751: color = 12'h000;
            1752: color = 12'h000;
            1753: color = 12'h000;
            1754: color = 12'h000;
            1755: color = 12'h000;
            1756: color = 12'h000;
            1757: color = 12'h000;
            1758: color = 12'h000;
            1759: color = 12'h000;
            1760: color = 12'h000;
            1761: color = 12'h000;
            1762: color = 12'h000;
            1763: color = 12'h000;
            1764: color = 12'h000;
            1765: color = 12'h000;
            1766: color = 12'h000;
            1767: color = 12'h000;
            1768: color = 12'h000;
            1769: color = 12'h000;
            1770: color = 12'h000;
            1771: color = 12'h000;
            1772: color = 12'h000;
            1773: color = 12'h000;
            1774: color = 12'h000;
            1775: color = 12'h000;
            1776: color = 12'h000;
            1777: color = 12'h000;
            1778: color = 12'h000;
            1779: color = 12'h000;
            1780: color = 12'h000;
            1781: color = 12'h000;
            1782: color = 12'h000;
            1783: color = 12'h000;
            1784: color = 12'h000;
            1785: color = 12'h000;
            1786: color = 12'h000;
            1787: color = 12'h000;
            1788: color = 12'h000;
            1789: color = 12'h000;
            1790: color = 12'h000;
            1791: color = 12'h000;
            1792: color = 12'h000;
            1793: color = 12'h000;
            1794: color = 12'h000;
            1795: color = 12'h000;
            1796: color = 12'h000;
            1797: color = 12'h000;
            1798: color = 12'h000;
            1799: color = 12'h000;
            1800: color = 12'h000;
            1801: color = 12'h000;
            1802: color = 12'h000;
            1803: color = 12'h000;
            1804: color = 12'h000;
            1805: color = 12'h000;
            1806: color = 12'h000;
            1807: color = 12'h000;
            1808: color = 12'h000;
            1809: color = 12'h000;
            1810: color = 12'h000;
            1811: color = 12'h000;
            1812: color = 12'h000;
            1813: color = 12'h000;
            1814: color = 12'h000;
            1815: color = 12'h000;
            1816: color = 12'h000;
            1817: color = 12'h000;
            1818: color = 12'h000;
            1819: color = 12'h000;
            1820: color = 12'h000;
            1821: color = 12'h000;
            1822: color = 12'h000;
            1823: color = 12'h000;
            1824: color = 12'h000;
            1825: color = 12'h000;
            1826: color = 12'h000;
            1827: color = 12'h000;
            1828: color = 12'h000;
            1829: color = 12'h000;
            1830: color = 12'h000;
            1831: color = 12'h000;
            1832: color = 12'h000;
            1833: color = 12'h000;
            1834: color = 12'h000;
            1835: color = 12'h000;
            1836: color = 12'h000;
            1837: color = 12'h000;
            1838: color = 12'h000;
            1839: color = 12'h000;
            1840: color = 12'h000;
            1841: color = 12'h000;
            1842: color = 12'h000;
            1843: color = 12'h000;
            1844: color = 12'h000;
            1845: color = 12'h000;
            1846: color = 12'h000;
            1847: color = 12'h000;
            1848: color = 12'h000;
            1849: color = 12'h000;
            1850: color = 12'h000;
            1851: color = 12'h000;
            1852: color = 12'h000;
            1853: color = 12'h000;
            1854: color = 12'h000;
            1855: color = 12'h000;
            1856: color = 12'h000;
            1857: color = 12'h000;
            1858: color = 12'h000;
            1859: color = 12'h000;
            1860: color = 12'h000;
            1861: color = 12'h000;
            1862: color = 12'h000;
            1863: color = 12'h000;
            1864: color = 12'h000;
            1865: color = 12'h000;
            1866: color = 12'h000;
            1867: color = 12'h000;
            1868: color = 12'h000;
            1869: color = 12'h000;
            1870: color = 12'h000;
            1871: color = 12'h000;
            1872: color = 12'h000;
            1873: color = 12'h000;
            1874: color = 12'h000;
            1875: color = 12'h000;
            1876: color = 12'h000;
            1877: color = 12'h000;
            1878: color = 12'h000;
            1879: color = 12'h000;
            1880: color = 12'h000;
            1881: color = 12'h000;
            1882: color = 12'h000;
            1883: color = 12'h000;
            1884: color = 12'h000;
            1885: color = 12'h000;
            1886: color = 12'h000;
            1887: color = 12'h000;
            1888: color = 12'h000;
            1889: color = 12'h000;
            1890: color = 12'h000;
            1891: color = 12'h000;
            1892: color = 12'h000;
            1893: color = 12'h000;
            1894: color = 12'h000;
            1895: color = 12'h000;
            1896: color = 12'h000;
            1897: color = 12'h000;
            1898: color = 12'h000;
            1899: color = 12'h000;
            1900: color = 12'h000;
            1901: color = 12'h000;
            1902: color = 12'h000;
            1903: color = 12'h000;
            1904: color = 12'h000;
            1905: color = 12'h000;
            1906: color = 12'h000;
            1907: color = 12'h000;
            1908: color = 12'h000;
            1909: color = 12'h000;
            1910: color = 12'h000;
            1911: color = 12'h000;
            1912: color = 12'h000;
            1913: color = 12'h000;
            1914: color = 12'h000;
            1915: color = 12'h000;
            1916: color = 12'h000;
            1917: color = 12'h000;
            1918: color = 12'h000;
            1919: color = 12'h000;
            1920: color = 12'h000;
            1921: color = 12'h000;
            1922: color = 12'h000;
            1923: color = 12'h000;
            1924: color = 12'h000;
            1925: color = 12'h000;
            1926: color = 12'h000;
            1927: color = 12'h000;
            1928: color = 12'h000;
            1929: color = 12'h000;
            1930: color = 12'h000;
            1931: color = 12'h000;
            1932: color = 12'h000;
            1933: color = 12'h000;
            1934: color = 12'h000;
            1935: color = 12'h000;
            1936: color = 12'h000;
            1937: color = 12'h000;
            1938: color = 12'h000;
            1939: color = 12'h000;
            1940: color = 12'h000;
            1941: color = 12'h000;
            1942: color = 12'h000;
            1943: color = 12'h000;
            1944: color = 12'h000;
            1945: color = 12'h000;
            1946: color = 12'h000;
            1947: color = 12'h000;
            1948: color = 12'h000;
            1949: color = 12'h000;
            1950: color = 12'h000;
            1951: color = 12'h000;
            1952: color = 12'h000;
            1953: color = 12'h000;
            1954: color = 12'h000;
            1955: color = 12'h000;
            1956: color = 12'h000;
            1957: color = 12'h000;
            1958: color = 12'h000;
            1959: color = 12'h000;
            1960: color = 12'h000;
            1961: color = 12'h000;
            1962: color = 12'h000;
            1963: color = 12'h000;
            1964: color = 12'h000;
            1965: color = 12'h000;
            1966: color = 12'h000;
            1967: color = 12'h000;
            1968: color = 12'h000;
            1969: color = 12'h000;
            1970: color = 12'h000;
            1971: color = 12'h000;
            1972: color = 12'h000;
            1973: color = 12'h000;
            1974: color = 12'h000;
            1975: color = 12'h000;
            1976: color = 12'h000;
            1977: color = 12'h000;
            1978: color = 12'h000;
            1979: color = 12'h000;
            1980: color = 12'h000;
            1981: color = 12'h000;
            1982: color = 12'h000;
            1983: color = 12'h000;
            1984: color = 12'h000;
            1985: color = 12'h000;
            1986: color = 12'h000;
            1987: color = 12'h000;
            1988: color = 12'h000;
            1989: color = 12'h000;
            1990: color = 12'h000;
            1991: color = 12'h000;
            1992: color = 12'h000;
            1993: color = 12'h000;
            1994: color = 12'h000;
            1995: color = 12'h000;
            1996: color = 12'h000;
            1997: color = 12'h000;
            1998: color = 12'h000;
            1999: color = 12'h000;
            2000: color = 12'h000;
            2001: color = 12'h000;
            2002: color = 12'h000;
            2003: color = 12'h000;
            2004: color = 12'h000;
            2005: color = 12'h000;
            2006: color = 12'h000;
            2007: color = 12'h000;
            2008: color = 12'h000;
            2009: color = 12'h000;
            2010: color = 12'h000;
            2011: color = 12'h000;
            2012: color = 12'h000;
            2013: color = 12'h000;
            2014: color = 12'h000;
            2015: color = 12'h000;
            2016: color = 12'h000;
            2017: color = 12'h000;
            2018: color = 12'h000;
            2019: color = 12'h000;
            2020: color = 12'h000;
            2021: color = 12'h000;
            2022: color = 12'h000;
            2023: color = 12'h000;
            2024: color = 12'h000;
            2025: color = 12'h000;
            2026: color = 12'h000;
            2027: color = 12'h000;
            2028: color = 12'h000;
            2029: color = 12'h000;
            2030: color = 12'h000;
            2031: color = 12'h000;
            2032: color = 12'h000;
            2033: color = 12'h000;
            2034: color = 12'h000;
            2035: color = 12'h000;
            2036: color = 12'h000;
            2037: color = 12'h000;
            2038: color = 12'h000;
            2039: color = 12'h000;
            2040: color = 12'h000;
            2041: color = 12'h000;
            2042: color = 12'h000;
            2043: color = 12'h000;
            2044: color = 12'h000;
            2045: color = 12'h000;
            2046: color = 12'h000;
            2047: color = 12'h000;
            2048: color = 12'h000;
            2049: color = 12'h000;
            2050: color = 12'h000;
            2051: color = 12'h000;
            2052: color = 12'h000;
            2053: color = 12'h000;
            2054: color = 12'h000;
            2055: color = 12'h000;
            2056: color = 12'h000;
            2057: color = 12'h000;
            2058: color = 12'h000;
            2059: color = 12'h000;
            2060: color = 12'h000;
            2061: color = 12'h000;
            2062: color = 12'h000;
            2063: color = 12'h000;
            2064: color = 12'h000;
            2065: color = 12'h000;
            2066: color = 12'h000;
            2067: color = 12'h000;
            2068: color = 12'h000;
            2069: color = 12'h000;
            2070: color = 12'h000;
            2071: color = 12'h000;
            2072: color = 12'h000;
            2073: color = 12'h000;
            2074: color = 12'h000;
            2075: color = 12'h000;
            2076: color = 12'h000;
            2077: color = 12'h000;
            2078: color = 12'h000;
            2079: color = 12'h000;
            2080: color = 12'h000;
            2081: color = 12'h000;
            2082: color = 12'h000;
            2083: color = 12'h000;
            2084: color = 12'h000;
            2085: color = 12'h000;
            2086: color = 12'h000;
            2087: color = 12'h000;
            2088: color = 12'h000;
            2089: color = 12'h000;
            2090: color = 12'h000;
            2091: color = 12'h000;
            2092: color = 12'h000;
            2093: color = 12'h000;
            2094: color = 12'h000;
            2095: color = 12'h000;
            2096: color = 12'h000;
            2097: color = 12'h000;
            2098: color = 12'h000;
            2099: color = 12'h000;
            2100: color = 12'h000;
            2101: color = 12'h000;
            2102: color = 12'h000;
            2103: color = 12'h000;
            2104: color = 12'h000;
            2105: color = 12'h000;
            2106: color = 12'h000;
            2107: color = 12'h000;
            2108: color = 12'h000;
            2109: color = 12'h000;
            2110: color = 12'h000;
            2111: color = 12'h000;
            2112: color = 12'h000;
            2113: color = 12'h000;
            2114: color = 12'h000;
            2115: color = 12'h000;
            2116: color = 12'h000;
            2117: color = 12'h000;
            2118: color = 12'h000;
            2119: color = 12'h000;
            2120: color = 12'h000;
            2121: color = 12'h000;
            2122: color = 12'h000;
            2123: color = 12'h000;
            2124: color = 12'h000;
            2125: color = 12'h000;
            2126: color = 12'h000;
            2127: color = 12'h000;
            2128: color = 12'h000;
            2129: color = 12'h000;
            2130: color = 12'h000;
            2131: color = 12'h000;
            2132: color = 12'h000;
            2133: color = 12'h000;
            2134: color = 12'h000;
            2135: color = 12'h000;
            2136: color = 12'h000;
            2137: color = 12'h000;
            2138: color = 12'h000;
            2139: color = 12'h000;
            2140: color = 12'h000;
            2141: color = 12'h000;
            2142: color = 12'h000;
            2143: color = 12'h000;
            2144: color = 12'h000;
            2145: color = 12'h000;
            2146: color = 12'h000;
            2147: color = 12'h000;
            2148: color = 12'h000;
            2149: color = 12'h000;
            2150: color = 12'h000;
            2151: color = 12'h000;
            2152: color = 12'h000;
            2153: color = 12'h000;
            2154: color = 12'h000;
            2155: color = 12'h000;
            2156: color = 12'h000;
            2157: color = 12'h000;
            2158: color = 12'h000;
            2159: color = 12'h000;
            2160: color = 12'h000;
            2161: color = 12'h000;
            2162: color = 12'h000;
            2163: color = 12'h000;
            2164: color = 12'h000;
            2165: color = 12'h000;
            2166: color = 12'h000;
            2167: color = 12'h000;
            2168: color = 12'h000;
            2169: color = 12'h000;
            2170: color = 12'h000;
            2171: color = 12'h000;
            2172: color = 12'h000;
            2173: color = 12'h000;
            2174: color = 12'h000;
            2175: color = 12'h000;
            2176: color = 12'h000;
            2177: color = 12'h000;
            2178: color = 12'h000;
            2179: color = 12'h000;
            2180: color = 12'h000;
            2181: color = 12'h000;
            2182: color = 12'h000;
            2183: color = 12'h000;
            2184: color = 12'h000;
            2185: color = 12'h000;
            2186: color = 12'h000;
            2187: color = 12'h000;
            2188: color = 12'h000;
            2189: color = 12'h000;
            2190: color = 12'h000;
            2191: color = 12'h000;
            2192: color = 12'h000;
            2193: color = 12'h000;
            2194: color = 12'h000;
            2195: color = 12'h000;
            2196: color = 12'h000;
            2197: color = 12'h000;
            2198: color = 12'h000;
            2199: color = 12'h000;
            2200: color = 12'h000;
            2201: color = 12'h000;
            2202: color = 12'h000;
            2203: color = 12'h000;
            2204: color = 12'h000;
            2205: color = 12'h000;
            2206: color = 12'h000;
            2207: color = 12'h000;
            2208: color = 12'h000;
            2209: color = 12'h000;
            2210: color = 12'h000;
            2211: color = 12'h000;
            2212: color = 12'h000;
            2213: color = 12'h000;
            2214: color = 12'h000;
            2215: color = 12'h000;
            2216: color = 12'h000;
            2217: color = 12'h000;
            2218: color = 12'h000;
            2219: color = 12'h000;
            2220: color = 12'h000;
            2221: color = 12'h000;
            2222: color = 12'h000;
            2223: color = 12'h000;
            2224: color = 12'h000;
            2225: color = 12'h000;
            2226: color = 12'h000;
            2227: color = 12'h000;
            2228: color = 12'h000;
            2229: color = 12'h000;
            2230: color = 12'h000;
            2231: color = 12'h000;
            2232: color = 12'h000;
            2233: color = 12'h000;
            2234: color = 12'h000;
            2235: color = 12'h000;
            2236: color = 12'h000;
            2237: color = 12'h000;
            2238: color = 12'h000;
            2239: color = 12'h000;
            2240: color = 12'h000;
            2241: color = 12'h000;
            2242: color = 12'h000;
            2243: color = 12'h000;
            2244: color = 12'h000;
            2245: color = 12'h000;
            2246: color = 12'h000;
            2247: color = 12'h000;
            2248: color = 12'h000;
            2249: color = 12'h000;
            2250: color = 12'h000;
            2251: color = 12'h000;
            2252: color = 12'h000;
            2253: color = 12'h000;
            2254: color = 12'h000;
            2255: color = 12'h000;
            2256: color = 12'h000;
            2257: color = 12'h000;
            2258: color = 12'h000;
            2259: color = 12'h000;
            2260: color = 12'h000;
            2261: color = 12'h000;
            2262: color = 12'h000;
            2263: color = 12'h000;
            2264: color = 12'h000;
            2265: color = 12'h000;
            2266: color = 12'h000;
            2267: color = 12'h000;
            2268: color = 12'h000;
            2269: color = 12'h000;
            2270: color = 12'h000;
            2271: color = 12'h000;
            2272: color = 12'h000;
            2273: color = 12'h000;
            2274: color = 12'h000;
            2275: color = 12'h000;
            2276: color = 12'h000;
            2277: color = 12'h000;
            2278: color = 12'h000;
            2279: color = 12'h000;
            2280: color = 12'h000;
            2281: color = 12'h000;
            2282: color = 12'h000;
            2283: color = 12'h000;
            2284: color = 12'h000;
            2285: color = 12'h000;
            2286: color = 12'h000;
            2287: color = 12'h000;
            2288: color = 12'h000;
            2289: color = 12'h000;
            2290: color = 12'h000;
            2291: color = 12'h000;
            2292: color = 12'h000;
            2293: color = 12'h000;
            2294: color = 12'h000;
            2295: color = 12'h000;
            2296: color = 12'h000;
            2297: color = 12'h000;
            2298: color = 12'h000;
            2299: color = 12'h000;
            2300: color = 12'h000;
            2301: color = 12'h000;
            2302: color = 12'h000;
            2303: color = 12'h000;
            2304: color = 12'h000;
            2305: color = 12'h000;
            2306: color = 12'h000;
            2307: color = 12'h000;
            2308: color = 12'h000;
            2309: color = 12'h000;
            2310: color = 12'h000;
            2311: color = 12'h000;
            2312: color = 12'h000;
            2313: color = 12'h000;
            2314: color = 12'h000;
            2315: color = 12'h000;
            2316: color = 12'h000;
            2317: color = 12'h000;
            2318: color = 12'h000;
            2319: color = 12'h000;
            2320: color = 12'h000;
            2321: color = 12'h000;
            2322: color = 12'h000;
            2323: color = 12'h000;
            2324: color = 12'h000;
            2325: color = 12'h000;
            2326: color = 12'h000;
            2327: color = 12'h000;
            2328: color = 12'h000;
            2329: color = 12'h000;
            2330: color = 12'h000;
            2331: color = 12'h000;
            2332: color = 12'h000;
            2333: color = 12'h000;
            2334: color = 12'h000;
            2335: color = 12'h000;
            2336: color = 12'h000;
            2337: color = 12'h000;
            2338: color = 12'h000;
            2339: color = 12'h000;
            2340: color = 12'h000;
            2341: color = 12'h000;
            2342: color = 12'h000;
            2343: color = 12'h000;
            2344: color = 12'h000;
            2345: color = 12'h000;
            2346: color = 12'h000;
            2347: color = 12'h000;
            2348: color = 12'h000;
            2349: color = 12'h000;
            2350: color = 12'h000;
            2351: color = 12'h000;
            2352: color = 12'h000;
            2353: color = 12'h000;
            2354: color = 12'h000;
            2355: color = 12'h000;
            2356: color = 12'h000;
            2357: color = 12'h000;
            2358: color = 12'h000;
            2359: color = 12'h000;
            2360: color = 12'h000;
            2361: color = 12'h000;
            2362: color = 12'h000;
            2363: color = 12'h000;
            2364: color = 12'h000;
            2365: color = 12'h000;
            2366: color = 12'h000;
            2367: color = 12'h000;
            2368: color = 12'h000;
            2369: color = 12'h000;
            2370: color = 12'h000;
            2371: color = 12'h000;
            2372: color = 12'h000;
            2373: color = 12'h000;
            2374: color = 12'h000;
            2375: color = 12'h000;
            2376: color = 12'h000;
            2377: color = 12'h000;
            2378: color = 12'h000;
            2379: color = 12'h000;
            2380: color = 12'h000;
            2381: color = 12'h000;
            2382: color = 12'h000;
            2383: color = 12'h000;
            2384: color = 12'h000;
            2385: color = 12'h000;
            2386: color = 12'h000;
            2387: color = 12'h000;
            2388: color = 12'h000;
            2389: color = 12'h000;
            2390: color = 12'h000;
            2391: color = 12'h000;
            2392: color = 12'h000;
            2393: color = 12'h000;
            2394: color = 12'h000;
            2395: color = 12'h000;
            2396: color = 12'h000;
            2397: color = 12'h000;
            2398: color = 12'h000;
            2399: color = 12'h000;
            2400: color = 12'h000;
            2401: color = 12'h000;
            2402: color = 12'h000;
            2403: color = 12'h000;
            2404: color = 12'h000;
            2405: color = 12'h000;
            2406: color = 12'h000;
            2407: color = 12'h000;
            2408: color = 12'h000;
            2409: color = 12'h000;
            2410: color = 12'h000;
            2411: color = 12'h000;
            2412: color = 12'h000;
            2413: color = 12'h000;
            2414: color = 12'h000;
            2415: color = 12'h000;
            2416: color = 12'h000;
            2417: color = 12'h000;
            2418: color = 12'h000;
            2419: color = 12'h000;
            2420: color = 12'h000;
            2421: color = 12'h000;
            2422: color = 12'h000;
            2423: color = 12'h000;
            2424: color = 12'h000;
            2425: color = 12'h000;
            2426: color = 12'h000;
            2427: color = 12'h000;
            2428: color = 12'h000;
            2429: color = 12'h000;
            2430: color = 12'h000;
            2431: color = 12'h000;
            2432: color = 12'h000;
            2433: color = 12'h000;
            2434: color = 12'h000;
            2435: color = 12'h000;
            2436: color = 12'h000;
            2437: color = 12'h000;
            2438: color = 12'h000;
            2439: color = 12'h000;
            2440: color = 12'h000;
            2441: color = 12'h000;
            2442: color = 12'h000;
            2443: color = 12'h000;
            2444: color = 12'h000;
            2445: color = 12'h000;
            2446: color = 12'h000;
            2447: color = 12'h000;
            2448: color = 12'h000;
            2449: color = 12'h000;
            2450: color = 12'h000;
            2451: color = 12'h000;
            2452: color = 12'h000;
            2453: color = 12'h000;
            2454: color = 12'h000;
            2455: color = 12'h000;
            2456: color = 12'h000;
            2457: color = 12'h000;
            2458: color = 12'h000;
            2459: color = 12'h000;
            2460: color = 12'h000;
            2461: color = 12'h000;
            2462: color = 12'h000;
            2463: color = 12'h000;
            2464: color = 12'h000;
            2465: color = 12'h000;
            2466: color = 12'h000;
            2467: color = 12'h000;
            2468: color = 12'h000;
            2469: color = 12'h000;
            2470: color = 12'h000;
            2471: color = 12'h000;
            2472: color = 12'h000;
            2473: color = 12'h000;
            2474: color = 12'h000;
            2475: color = 12'h000;
            2476: color = 12'h000;
            2477: color = 12'h000;
            2478: color = 12'h000;
            2479: color = 12'h000;
            2480: color = 12'h000;
            2481: color = 12'h000;
            2482: color = 12'h000;
            2483: color = 12'h000;
            2484: color = 12'h000;
            2485: color = 12'h000;
            2486: color = 12'h000;
            2487: color = 12'h000;
            2488: color = 12'h000;
            2489: color = 12'h000;
            2490: color = 12'h000;
            2491: color = 12'h000;
            2492: color = 12'h000;
            2493: color = 12'h000;
            2494: color = 12'h000;
            2495: color = 12'h000;
            2496: color = 12'h000;
            2497: color = 12'h000;
            2498: color = 12'h000;
            2499: color = 12'h000;
            2500: color = 12'h000;
            2501: color = 12'h000;
            2502: color = 12'h000;
            2503: color = 12'h000;
            2504: color = 12'h000;
            2505: color = 12'h000;
            2506: color = 12'h000;
            2507: color = 12'h000;
            2508: color = 12'h000;
            2509: color = 12'h000;
            2510: color = 12'h000;
            2511: color = 12'h000;
            2512: color = 12'h000;
            2513: color = 12'h000;
            2514: color = 12'h000;
            2515: color = 12'h000;
            2516: color = 12'h000;
            2517: color = 12'h000;
            2518: color = 12'h000;
            2519: color = 12'h000;
            2520: color = 12'h000;
            2521: color = 12'h000;
            2522: color = 12'h000;
            2523: color = 12'h000;
            2524: color = 12'h000;
            2525: color = 12'h000;
            2526: color = 12'h000;
            2527: color = 12'h000;
            2528: color = 12'h000;
            2529: color = 12'h000;
            2530: color = 12'h000;
            2531: color = 12'h000;
            2532: color = 12'h000;
            2533: color = 12'h000;
            2534: color = 12'h000;
            2535: color = 12'h000;
            2536: color = 12'h000;
            2537: color = 12'h000;
            2538: color = 12'h000;
            2539: color = 12'h000;
            2540: color = 12'h000;
            2541: color = 12'h000;
            2542: color = 12'h000;
            2543: color = 12'h000;
            2544: color = 12'h000;
            2545: color = 12'h000;
            2546: color = 12'h000;
            2547: color = 12'h000;
            2548: color = 12'h000;
            2549: color = 12'h000;
            2550: color = 12'h000;
            2551: color = 12'h000;
            2552: color = 12'h000;
            2553: color = 12'h000;
            2554: color = 12'h000;
            2555: color = 12'h000;
            2556: color = 12'h000;
            2557: color = 12'h000;
            2558: color = 12'h000;
            2559: color = 12'h000;
            2560: color = 12'h000;
            2561: color = 12'h000;
            2562: color = 12'h000;
            2563: color = 12'h000;
            2564: color = 12'h000;
            2565: color = 12'h000;
            2566: color = 12'h000;
            2567: color = 12'h000;
            2568: color = 12'h000;
            2569: color = 12'h000;
            2570: color = 12'h000;
            2571: color = 12'h000;
            2572: color = 12'h000;
            2573: color = 12'h000;
            2574: color = 12'h000;
            2575: color = 12'h000;
            2576: color = 12'h000;
            2577: color = 12'h000;
            2578: color = 12'h000;
            2579: color = 12'h000;
            2580: color = 12'h000;
            2581: color = 12'h000;
            2582: color = 12'h000;
            2583: color = 12'h000;
            2584: color = 12'h000;
            2585: color = 12'h000;
            2586: color = 12'h000;
            2587: color = 12'h000;
            2588: color = 12'h000;
            2589: color = 12'h000;
            2590: color = 12'h000;
            2591: color = 12'h000;
            2592: color = 12'h000;
            2593: color = 12'h000;
            2594: color = 12'h000;
            2595: color = 12'h000;
            2596: color = 12'h000;
            2597: color = 12'h000;
            2598: color = 12'h000;
            2599: color = 12'h000;
            2600: color = 12'h000;
            2601: color = 12'h000;
            2602: color = 12'h000;
            2603: color = 12'h000;
            2604: color = 12'h000;
            2605: color = 12'h000;
            2606: color = 12'h000;
            2607: color = 12'h000;
            2608: color = 12'h000;
            2609: color = 12'h000;
            2610: color = 12'h000;
            2611: color = 12'h000;
            2612: color = 12'h000;
            2613: color = 12'h000;
            2614: color = 12'h000;
            2615: color = 12'h000;
            2616: color = 12'h000;
            2617: color = 12'h000;
            2618: color = 12'h000;
            2619: color = 12'h000;
            2620: color = 12'h000;
            2621: color = 12'h000;
            2622: color = 12'h000;
            2623: color = 12'h000;
            2624: color = 12'h000;
            2625: color = 12'h000;
            2626: color = 12'h000;
            2627: color = 12'h000;
            2628: color = 12'h000;
            2629: color = 12'h000;
            2630: color = 12'h000;
            2631: color = 12'h000;
            2632: color = 12'h000;
            2633: color = 12'h000;
            2634: color = 12'h000;
            2635: color = 12'h000;
            2636: color = 12'h000;
            2637: color = 12'h000;
            2638: color = 12'h000;
            2639: color = 12'h000;
            2640: color = 12'h000;
            2641: color = 12'h000;
            2642: color = 12'h000;
            2643: color = 12'h000;
            2644: color = 12'h000;
            2645: color = 12'h000;
            2646: color = 12'h000;
            2647: color = 12'h000;
            2648: color = 12'h000;
            2649: color = 12'h000;
            2650: color = 12'h000;
            2651: color = 12'h000;
            2652: color = 12'h000;
            2653: color = 12'h000;
            2654: color = 12'h000;
            2655: color = 12'h000;
            2656: color = 12'h000;
            2657: color = 12'h000;
            2658: color = 12'h000;
            2659: color = 12'h000;
            2660: color = 12'h000;
            2661: color = 12'h000;
            2662: color = 12'h000;
            2663: color = 12'h000;
            2664: color = 12'h000;
            2665: color = 12'h000;
            2666: color = 12'h000;
            2667: color = 12'h000;
            2668: color = 12'h000;
            2669: color = 12'h000;
            2670: color = 12'h000;
            2671: color = 12'h000;
            2672: color = 12'h000;
            2673: color = 12'h000;
            2674: color = 12'h000;
            2675: color = 12'h000;
            2676: color = 12'h000;
            2677: color = 12'h000;
            2678: color = 12'h000;
            2679: color = 12'h000;
            2680: color = 12'h000;
            2681: color = 12'h000;
            2682: color = 12'h000;
            2683: color = 12'h000;
            2684: color = 12'h000;
            2685: color = 12'h000;
            2686: color = 12'h000;
            2687: color = 12'h000;
            2688: color = 12'h000;
            2689: color = 12'h000;
            2690: color = 12'h000;
            2691: color = 12'h000;
            2692: color = 12'h000;
            2693: color = 12'h000;
            2694: color = 12'h000;
            2695: color = 12'h000;
            2696: color = 12'h000;
            2697: color = 12'h000;
            2698: color = 12'h000;
            2699: color = 12'h000;
            2700: color = 12'h000;
            2701: color = 12'h000;
            2702: color = 12'h000;
            2703: color = 12'h000;
            2704: color = 12'h000;
            2705: color = 12'h000;
            2706: color = 12'h000;
            2707: color = 12'h000;
            2708: color = 12'h000;
            2709: color = 12'h000;
            2710: color = 12'h000;
            2711: color = 12'h000;
            2712: color = 12'h000;
            2713: color = 12'h000;
            2714: color = 12'h000;
            2715: color = 12'h000;
            2716: color = 12'h000;
            2717: color = 12'h000;
            2718: color = 12'h000;
            2719: color = 12'h000;
            2720: color = 12'h000;
            2721: color = 12'h000;
            2722: color = 12'h000;
            2723: color = 12'h000;
            2724: color = 12'h000;
            2725: color = 12'h000;
            2726: color = 12'h000;
            2727: color = 12'h000;
            2728: color = 12'h000;
            2729: color = 12'h000;
            2730: color = 12'h000;
            2731: color = 12'h000;
            2732: color = 12'h000;
            2733: color = 12'h000;
            2734: color = 12'h000;
            2735: color = 12'h000;
            2736: color = 12'h000;
            2737: color = 12'h000;
            2738: color = 12'h000;
            2739: color = 12'h000;
            2740: color = 12'h000;
            2741: color = 12'h000;
            2742: color = 12'h000;
            2743: color = 12'h000;
            2744: color = 12'h000;
            2745: color = 12'h000;
            2746: color = 12'h000;
            2747: color = 12'h000;
            2748: color = 12'h000;
            2749: color = 12'h000;
            2750: color = 12'h000;
            2751: color = 12'h000;
            2752: color = 12'h000;
            2753: color = 12'h000;
            2754: color = 12'h000;
            2755: color = 12'h000;
            2756: color = 12'h000;
            2757: color = 12'h000;
            2758: color = 12'h000;
            2759: color = 12'h000;
            2760: color = 12'h000;
            2761: color = 12'h000;
            2762: color = 12'h000;
            2763: color = 12'h000;
            2764: color = 12'h000;
            2765: color = 12'h000;
            2766: color = 12'h000;
            2767: color = 12'h000;
            2768: color = 12'h000;
            2769: color = 12'h000;
            2770: color = 12'h000;
            2771: color = 12'h000;
            2772: color = 12'h000;
            2773: color = 12'h000;
            2774: color = 12'h000;
            2775: color = 12'h000;
            2776: color = 12'h000;
            2777: color = 12'h000;
            2778: color = 12'h000;
            2779: color = 12'h000;
            2780: color = 12'h000;
            2781: color = 12'h000;
            2782: color = 12'h000;
            2783: color = 12'h000;
            2784: color = 12'h000;
            2785: color = 12'h000;
            2786: color = 12'h000;
            2787: color = 12'h000;
            2788: color = 12'h000;
            2789: color = 12'h000;
            2790: color = 12'h000;
            2791: color = 12'h000;
            2792: color = 12'h000;
            2793: color = 12'h000;
            2794: color = 12'h000;
            2795: color = 12'h000;
            2796: color = 12'h000;
            2797: color = 12'h000;
            2798: color = 12'h000;
            2799: color = 12'h000;
            2800: color = 12'h000;
            2801: color = 12'h000;
            2802: color = 12'h000;
            2803: color = 12'h000;
            2804: color = 12'h000;
            2805: color = 12'h000;
            2806: color = 12'h000;
            2807: color = 12'h000;
            2808: color = 12'h000;
            2809: color = 12'h000;
            2810: color = 12'h000;
            2811: color = 12'h000;
            2812: color = 12'h000;
            2813: color = 12'h000;
            2814: color = 12'h000;
            2815: color = 12'h000;
            2816: color = 12'h000;
            2817: color = 12'h000;
            2818: color = 12'h000;
            2819: color = 12'h000;
            2820: color = 12'h000;
            2821: color = 12'h000;
            2822: color = 12'h000;
            2823: color = 12'h000;
            2824: color = 12'h000;
            2825: color = 12'h000;
            2826: color = 12'h000;
            2827: color = 12'h000;
            2828: color = 12'h000;
            2829: color = 12'h000;
            2830: color = 12'h000;
            2831: color = 12'h000;
            2832: color = 12'h000;
            2833: color = 12'h000;
            2834: color = 12'h000;
            2835: color = 12'h000;
            2836: color = 12'h000;
            2837: color = 12'h000;
            2838: color = 12'h000;
            2839: color = 12'h000;
            2840: color = 12'h000;
            2841: color = 12'h000;
            2842: color = 12'h000;
            2843: color = 12'h000;
            2844: color = 12'h000;
            2845: color = 12'h000;
            2846: color = 12'h000;
            2847: color = 12'h000;
            2848: color = 12'h000;
            2849: color = 12'h000;
            2850: color = 12'h000;
            2851: color = 12'h000;
            2852: color = 12'h000;
            2853: color = 12'h000;
            2854: color = 12'h000;
            2855: color = 12'h000;
            2856: color = 12'h000;
            2857: color = 12'h000;
            2858: color = 12'h000;
            2859: color = 12'h000;
            2860: color = 12'h000;
            2861: color = 12'h000;
            2862: color = 12'h000;
            2863: color = 12'h000;
            2864: color = 12'h000;
            2865: color = 12'h000;
            2866: color = 12'h000;
            2867: color = 12'h000;
            2868: color = 12'h000;
            2869: color = 12'h000;
            2870: color = 12'h000;
            2871: color = 12'h000;
            2872: color = 12'h000;
            2873: color = 12'h000;
            2874: color = 12'h000;
            2875: color = 12'h000;
            2876: color = 12'h000;
            2877: color = 12'h000;
            2878: color = 12'h000;
            2879: color = 12'h000;
            2880: color = 12'h000;
            2881: color = 12'h000;
            2882: color = 12'h000;
            2883: color = 12'h000;
            2884: color = 12'h000;
            2885: color = 12'h000;
            2886: color = 12'h000;
            2887: color = 12'h000;
            2888: color = 12'h000;
            2889: color = 12'h000;
            2890: color = 12'h000;
            2891: color = 12'h000;
            2892: color = 12'h000;
            2893: color = 12'h000;
            2894: color = 12'h000;
            2895: color = 12'h000;
            2896: color = 12'h000;
            2897: color = 12'h000;
            2898: color = 12'h000;
            2899: color = 12'h000;
            2900: color = 12'h000;
            2901: color = 12'h000;
            2902: color = 12'h000;
            2903: color = 12'h000;
            2904: color = 12'h000;
            2905: color = 12'h000;
            2906: color = 12'h000;
            2907: color = 12'h000;
            2908: color = 12'h000;
            2909: color = 12'h000;
            2910: color = 12'h000;
            2911: color = 12'h000;
            2912: color = 12'h000;
            2913: color = 12'h000;
            2914: color = 12'h000;
            2915: color = 12'h000;
            2916: color = 12'h000;
            2917: color = 12'h000;
            2918: color = 12'h000;
            2919: color = 12'h000;
            2920: color = 12'h000;
            2921: color = 12'h000;
            2922: color = 12'h000;
            2923: color = 12'h000;
            2924: color = 12'h000;
            2925: color = 12'h000;
            2926: color = 12'h000;
            2927: color = 12'h000;
            2928: color = 12'h000;
            2929: color = 12'h000;
            2930: color = 12'h000;
            2931: color = 12'h000;
            2932: color = 12'h000;
            2933: color = 12'h000;
            2934: color = 12'h000;
            2935: color = 12'h000;
            2936: color = 12'h000;
            2937: color = 12'h000;
            2938: color = 12'h000;
            2939: color = 12'h000;
            2940: color = 12'h000;
            2941: color = 12'h000;
            2942: color = 12'h000;
            2943: color = 12'h000;
            2944: color = 12'h000;
            2945: color = 12'h000;
            2946: color = 12'h000;
            2947: color = 12'h000;
            2948: color = 12'h000;
            2949: color = 12'h000;
            2950: color = 12'h000;
            2951: color = 12'h000;
            2952: color = 12'h000;
            2953: color = 12'h000;
            2954: color = 12'h000;
            2955: color = 12'h000;
            2956: color = 12'h000;
            2957: color = 12'h000;
            2958: color = 12'h000;
            2959: color = 12'h000;
            2960: color = 12'h000;
            2961: color = 12'h000;
            2962: color = 12'h000;
            2963: color = 12'h000;
            2964: color = 12'h000;
            2965: color = 12'h000;
            2966: color = 12'h000;
            2967: color = 12'h000;
            2968: color = 12'h000;
            2969: color = 12'h000;
            2970: color = 12'h000;
            2971: color = 12'h000;
            2972: color = 12'h000;
            2973: color = 12'h000;
            2974: color = 12'h000;
            2975: color = 12'h000;
            2976: color = 12'h000;
            2977: color = 12'h000;
            2978: color = 12'h000;
            2979: color = 12'h000;
            2980: color = 12'h000;
            2981: color = 12'h000;
            2982: color = 12'h000;
            2983: color = 12'h000;
            2984: color = 12'h000;
            2985: color = 12'h000;
            2986: color = 12'h000;
            2987: color = 12'h000;
            2988: color = 12'h000;
            2989: color = 12'h000;
            2990: color = 12'h000;
            2991: color = 12'h000;
            2992: color = 12'h000;
            2993: color = 12'h000;
            2994: color = 12'h000;
            2995: color = 12'h000;
            2996: color = 12'h000;
            2997: color = 12'h000;
            2998: color = 12'h000;
            2999: color = 12'h000;
            3000: color = 12'h000;
            3001: color = 12'h000;
            3002: color = 12'h000;
            3003: color = 12'h000;
            3004: color = 12'h000;
            3005: color = 12'h000;
            3006: color = 12'h000;
            3007: color = 12'h000;
            3008: color = 12'h000;
            3009: color = 12'h000;
            3010: color = 12'h000;
            3011: color = 12'h000;
            3012: color = 12'h000;
            3013: color = 12'h000;
            3014: color = 12'h000;
            3015: color = 12'h000;
            3016: color = 12'h000;
            3017: color = 12'h000;
            3018: color = 12'h000;
            3019: color = 12'h000;
            3020: color = 12'h000;
            3021: color = 12'h000;
            3022: color = 12'h000;
            3023: color = 12'h000;
            3024: color = 12'h000;
            3025: color = 12'h000;
            3026: color = 12'h000;
            3027: color = 12'h000;
            3028: color = 12'h000;
            3029: color = 12'h000;
            3030: color = 12'h000;
            3031: color = 12'h000;
            3032: color = 12'h000;
            3033: color = 12'h000;
            3034: color = 12'h000;
            3035: color = 12'h000;
            3036: color = 12'h000;
            3037: color = 12'h000;
            3038: color = 12'h000;
            3039: color = 12'h000;
            3040: color = 12'h000;
            3041: color = 12'h000;
            3042: color = 12'h000;
            3043: color = 12'h000;
            3044: color = 12'h000;
            3045: color = 12'h000;
            3046: color = 12'h000;
            3047: color = 12'h000;
            3048: color = 12'h000;
            3049: color = 12'h000;
            3050: color = 12'h000;
            3051: color = 12'h000;
            3052: color = 12'h000;
            3053: color = 12'h000;
            3054: color = 12'h000;
            3055: color = 12'h000;
            3056: color = 12'h000;
            3057: color = 12'h000;
            3058: color = 12'h000;
            3059: color = 12'h000;
            3060: color = 12'h000;
            3061: color = 12'h000;
            3062: color = 12'h000;
            3063: color = 12'h000;
            3064: color = 12'h000;
            3065: color = 12'h000;
            3066: color = 12'h000;
            3067: color = 12'h000;
            3068: color = 12'h000;
            3069: color = 12'h000;
            3070: color = 12'h000;
            3071: color = 12'h000;
            3072: color = 12'h000;
            3073: color = 12'h000;
            3074: color = 12'h000;
            3075: color = 12'h000;
            3076: color = 12'h000;
            3077: color = 12'h000;
            3078: color = 12'h000;
            3079: color = 12'h000;
            3080: color = 12'h000;
            3081: color = 12'h000;
            3082: color = 12'h000;
            3083: color = 12'h000;
            3084: color = 12'h000;
            3085: color = 12'h000;
            3086: color = 12'h000;
            3087: color = 12'h000;
            3088: color = 12'h000;
            3089: color = 12'h000;
            3090: color = 12'h000;
            3091: color = 12'h000;
            3092: color = 12'h000;
            3093: color = 12'h000;
            3094: color = 12'h000;
            3095: color = 12'h000;
            3096: color = 12'h000;
            3097: color = 12'h000;
            3098: color = 12'h000;
            3099: color = 12'h000;
            3100: color = 12'h000;
            3101: color = 12'h000;
            3102: color = 12'h000;
            3103: color = 12'h000;
            3104: color = 12'h000;
            3105: color = 12'h000;
            3106: color = 12'h000;
            3107: color = 12'h000;
            3108: color = 12'h000;
            3109: color = 12'h000;
            3110: color = 12'h000;
            3111: color = 12'h000;
            3112: color = 12'h000;
            3113: color = 12'h000;
            3114: color = 12'h000;
            3115: color = 12'h000;
            3116: color = 12'h000;
            3117: color = 12'h000;
            3118: color = 12'h000;
            3119: color = 12'h000;
            3120: color = 12'h000;
            3121: color = 12'h000;
            3122: color = 12'h000;
            3123: color = 12'h000;
            3124: color = 12'h000;
            3125: color = 12'h000;
            3126: color = 12'h000;
            3127: color = 12'h000;
            3128: color = 12'h000;
            3129: color = 12'h000;
            3130: color = 12'h000;
            3131: color = 12'h000;
            3132: color = 12'h000;
            3133: color = 12'h000;
            3134: color = 12'h000;
            3135: color = 12'h000;
            3136: color = 12'h000;
            3137: color = 12'h000;
            3138: color = 12'h000;
            3139: color = 12'h000;
            3140: color = 12'h000;
            3141: color = 12'h000;
            3142: color = 12'h000;
            3143: color = 12'h000;
            3144: color = 12'h000;
            3145: color = 12'h000;
            3146: color = 12'h000;
            3147: color = 12'h000;
            3148: color = 12'h000;
            3149: color = 12'h000;
            3150: color = 12'h000;
            3151: color = 12'h000;
            3152: color = 12'h000;
            3153: color = 12'h000;
            3154: color = 12'h000;
            3155: color = 12'h000;
            3156: color = 12'h000;
            3157: color = 12'h000;
            3158: color = 12'h000;
            3159: color = 12'h000;
            3160: color = 12'h000;
            3161: color = 12'h000;
            3162: color = 12'h000;
            3163: color = 12'h000;
            3164: color = 12'h000;
            3165: color = 12'h000;
            3166: color = 12'h000;
            3167: color = 12'h000;
            3168: color = 12'h000;
            3169: color = 12'h000;
            3170: color = 12'h000;
            3171: color = 12'h000;
            3172: color = 12'h000;
            3173: color = 12'h000;
            3174: color = 12'h000;
            3175: color = 12'h000;
            3176: color = 12'h000;
            3177: color = 12'h000;
            3178: color = 12'h000;
            3179: color = 12'h000;
            3180: color = 12'h000;
            3181: color = 12'h000;
            3182: color = 12'h000;
            3183: color = 12'h000;
            3184: color = 12'h000;
            3185: color = 12'h000;
            3186: color = 12'h000;
            3187: color = 12'h000;
            3188: color = 12'h000;
            3189: color = 12'h000;
            3190: color = 12'h000;
            3191: color = 12'h000;
            3192: color = 12'h000;
            3193: color = 12'h000;
            3194: color = 12'h000;
            3195: color = 12'h000;
            3196: color = 12'h000;
            3197: color = 12'h000;
            3198: color = 12'h000;
            3199: color = 12'h000;
            3200: color = 12'h000;
            3201: color = 12'h000;
            3202: color = 12'h000;
            3203: color = 12'h000;
            3204: color = 12'h000;
            3205: color = 12'h000;
            3206: color = 12'h000;
            3207: color = 12'h000;
            3208: color = 12'h000;
            3209: color = 12'h000;
            3210: color = 12'h000;
            3211: color = 12'h000;
            3212: color = 12'h000;
            3213: color = 12'h000;
            3214: color = 12'h000;
            3215: color = 12'h000;
            3216: color = 12'h000;
            3217: color = 12'h000;
            3218: color = 12'h000;
            3219: color = 12'h000;
            3220: color = 12'h000;
            3221: color = 12'h000;
            3222: color = 12'h000;
            3223: color = 12'h000;
            3224: color = 12'h000;
            3225: color = 12'h000;
            3226: color = 12'h000;
            3227: color = 12'h000;
            3228: color = 12'h000;
            3229: color = 12'h000;
            3230: color = 12'h000;
            3231: color = 12'h000;
            3232: color = 12'h000;
            3233: color = 12'h000;
            3234: color = 12'h000;
            3235: color = 12'h000;
            3236: color = 12'h000;
            3237: color = 12'h000;
            3238: color = 12'h000;
            3239: color = 12'h000;
            3240: color = 12'h000;
            3241: color = 12'h000;
            3242: color = 12'h000;
            3243: color = 12'h000;
            3244: color = 12'h000;
            3245: color = 12'h000;
            3246: color = 12'h000;
            3247: color = 12'h000;
            3248: color = 12'h000;
            3249: color = 12'h000;
            3250: color = 12'h000;
            3251: color = 12'h000;
            3252: color = 12'h000;
            3253: color = 12'h000;
            3254: color = 12'h000;
            3255: color = 12'h000;
            3256: color = 12'h000;
            3257: color = 12'h000;
            3258: color = 12'h000;
            3259: color = 12'h000;
            3260: color = 12'h000;
            3261: color = 12'h000;
            3262: color = 12'h000;
            3263: color = 12'h000;
            3264: color = 12'h000;
            3265: color = 12'h000;
            3266: color = 12'h000;
            3267: color = 12'h000;
            3268: color = 12'h000;
            3269: color = 12'h000;
            3270: color = 12'h000;
            3271: color = 12'h000;
            3272: color = 12'h000;
            3273: color = 12'h000;
            3274: color = 12'h000;
            3275: color = 12'h000;
            3276: color = 12'h000;
            3277: color = 12'h000;
            3278: color = 12'h000;
            3279: color = 12'h000;
            3280: color = 12'h000;
            3281: color = 12'h000;
            3282: color = 12'h000;
            3283: color = 12'h000;
            3284: color = 12'h000;
            3285: color = 12'h000;
            3286: color = 12'h000;
            3287: color = 12'h000;
            3288: color = 12'h000;
            3289: color = 12'h000;
            3290: color = 12'h000;
            3291: color = 12'h000;
            3292: color = 12'h000;
            3293: color = 12'h000;
            3294: color = 12'h000;
            3295: color = 12'h000;
            3296: color = 12'h000;
            3297: color = 12'h000;
            3298: color = 12'h000;
            3299: color = 12'h000;
            3300: color = 12'h000;
            3301: color = 12'h000;
            3302: color = 12'h000;
            3303: color = 12'h000;
            3304: color = 12'h000;
            3305: color = 12'h000;
            3306: color = 12'h000;
            3307: color = 12'h000;
            3308: color = 12'h000;
            3309: color = 12'h000;
            3310: color = 12'h000;
            3311: color = 12'h000;
            3312: color = 12'h000;
            3313: color = 12'h000;
            3314: color = 12'h000;
            3315: color = 12'h000;
            3316: color = 12'h000;
            3317: color = 12'h000;
            3318: color = 12'h000;
            3319: color = 12'h000;
            3320: color = 12'h000;
            3321: color = 12'h000;
            3322: color = 12'h000;
            3323: color = 12'h000;
            3324: color = 12'h000;
            3325: color = 12'h000;
            3326: color = 12'h000;
            3327: color = 12'h000;
            3328: color = 12'h000;
            3329: color = 12'h000;
            3330: color = 12'h000;
            3331: color = 12'h000;
            3332: color = 12'h000;
            3333: color = 12'h000;
            3334: color = 12'h000;
            3335: color = 12'h000;
            3336: color = 12'h000;
            3337: color = 12'h000;
            3338: color = 12'h000;
            3339: color = 12'h000;
            3340: color = 12'h000;
            3341: color = 12'h000;
            3342: color = 12'h000;
            3343: color = 12'h000;
            3344: color = 12'h000;
            3345: color = 12'h000;
            3346: color = 12'h000;
            3347: color = 12'h000;
            3348: color = 12'h000;
            3349: color = 12'h000;
            3350: color = 12'h000;
            3351: color = 12'h000;
            3352: color = 12'h000;
            3353: color = 12'h000;
            3354: color = 12'h000;
            3355: color = 12'h000;
            3356: color = 12'h000;
            3357: color = 12'h000;
            3358: color = 12'h000;
            3359: color = 12'h000;
            3360: color = 12'h000;
            3361: color = 12'h000;
            3362: color = 12'h000;
            3363: color = 12'h000;
            3364: color = 12'h000;
            3365: color = 12'h000;
            3366: color = 12'h000;
            3367: color = 12'h000;
            3368: color = 12'h000;
            3369: color = 12'h000;
            3370: color = 12'h000;
            3371: color = 12'h000;
            3372: color = 12'h000;
            3373: color = 12'h000;
            3374: color = 12'h000;
            3375: color = 12'h000;
            3376: color = 12'h000;
            3377: color = 12'h000;
            3378: color = 12'h000;
            3379: color = 12'h000;
            3380: color = 12'h000;
            3381: color = 12'h000;
            3382: color = 12'h000;
            3383: color = 12'h000;
            3384: color = 12'h000;
            3385: color = 12'h000;
            3386: color = 12'h000;
            3387: color = 12'h000;
            3388: color = 12'h000;
            3389: color = 12'h000;
            3390: color = 12'h000;
            3391: color = 12'h000;
            3392: color = 12'h000;
            3393: color = 12'h000;
            3394: color = 12'h000;
            3395: color = 12'h000;
            3396: color = 12'h000;
            3397: color = 12'h000;
            3398: color = 12'h000;
            3399: color = 12'h000;
            3400: color = 12'h000;
            3401: color = 12'h000;
            3402: color = 12'h000;
            3403: color = 12'h000;
            3404: color = 12'h000;
            3405: color = 12'h000;
            3406: color = 12'h000;
            3407: color = 12'h000;
            3408: color = 12'h000;
            3409: color = 12'h000;
            3410: color = 12'h000;
            3411: color = 12'h000;
            3412: color = 12'h000;
            3413: color = 12'h000;
            3414: color = 12'h000;
            3415: color = 12'h000;
            3416: color = 12'h000;
            3417: color = 12'h000;
            3418: color = 12'h000;
            3419: color = 12'h000;
            3420: color = 12'h000;
            3421: color = 12'h000;
            3422: color = 12'h000;
            3423: color = 12'h000;
            3424: color = 12'h000;
            3425: color = 12'h000;
            3426: color = 12'h000;
            3427: color = 12'h000;
            3428: color = 12'h000;
            3429: color = 12'h000;
            3430: color = 12'h000;
            3431: color = 12'h000;
            3432: color = 12'h000;
            3433: color = 12'h000;
            3434: color = 12'h000;
            3435: color = 12'h000;
            3436: color = 12'h000;
            3437: color = 12'h000;
            3438: color = 12'h000;
            3439: color = 12'h000;
            3440: color = 12'h000;
            3441: color = 12'h000;
            3442: color = 12'h000;
            3443: color = 12'h000;
            3444: color = 12'h000;
            3445: color = 12'h000;
            3446: color = 12'h000;
            3447: color = 12'h000;
            3448: color = 12'h000;
            3449: color = 12'h000;
            3450: color = 12'h000;
            3451: color = 12'h000;
            3452: color = 12'h000;
            3453: color = 12'h000;
            3454: color = 12'h000;
            3455: color = 12'h000;
            3456: color = 12'h000;
            3457: color = 12'h000;
            3458: color = 12'h000;
            3459: color = 12'h000;
            3460: color = 12'h000;
            3461: color = 12'h000;
            3462: color = 12'h000;
            3463: color = 12'h000;
            3464: color = 12'h000;
            3465: color = 12'h000;
            3466: color = 12'h000;
            3467: color = 12'h000;
            3468: color = 12'h000;
            3469: color = 12'h000;
            3470: color = 12'h000;
            3471: color = 12'h000;
            3472: color = 12'h000;
            3473: color = 12'h000;
            3474: color = 12'h000;
            3475: color = 12'h000;
            3476: color = 12'h000;
            3477: color = 12'h000;
            3478: color = 12'h000;
            3479: color = 12'h000;
            3480: color = 12'h000;
            3481: color = 12'h000;
            3482: color = 12'h000;
            3483: color = 12'h000;
            3484: color = 12'h000;
            3485: color = 12'h000;
            3486: color = 12'h000;
            3487: color = 12'h000;
            3488: color = 12'h000;
            3489: color = 12'h000;
            3490: color = 12'h000;
            3491: color = 12'h000;
            3492: color = 12'h000;
            3493: color = 12'h000;
            3494: color = 12'h000;
            3495: color = 12'h000;
            3496: color = 12'h000;
            3497: color = 12'h000;
            3498: color = 12'h000;
            3499: color = 12'h000;
            3500: color = 12'h000;
            3501: color = 12'h000;
            3502: color = 12'h000;
            3503: color = 12'h000;
            3504: color = 12'h000;
            3505: color = 12'h000;
            3506: color = 12'h000;
            3507: color = 12'h000;
            3508: color = 12'h000;
            3509: color = 12'h000;
            3510: color = 12'h000;
            3511: color = 12'h000;
            3512: color = 12'h000;
            3513: color = 12'h000;
            3514: color = 12'h000;
            3515: color = 12'h000;
            3516: color = 12'h000;
            3517: color = 12'h000;
            3518: color = 12'h000;
            3519: color = 12'h000;
            3520: color = 12'h000;
            3521: color = 12'h000;
            3522: color = 12'h000;
            3523: color = 12'h000;
            3524: color = 12'h000;
            3525: color = 12'h000;
            3526: color = 12'h000;
            3527: color = 12'h000;
            3528: color = 12'h000;
            3529: color = 12'h000;
            3530: color = 12'h000;
            3531: color = 12'h000;
            3532: color = 12'h000;
            3533: color = 12'h000;
            3534: color = 12'h000;
            3535: color = 12'h000;
            3536: color = 12'h000;
            3537: color = 12'h000;
            3538: color = 12'h000;
            3539: color = 12'h000;
            3540: color = 12'h000;
            3541: color = 12'h000;
            3542: color = 12'h000;
            3543: color = 12'h000;
            3544: color = 12'h000;
            3545: color = 12'h000;
            3546: color = 12'h000;
            3547: color = 12'h000;
            3548: color = 12'h000;
            3549: color = 12'h000;
            3550: color = 12'h000;
            3551: color = 12'h000;
            3552: color = 12'h000;
            3553: color = 12'h000;
            3554: color = 12'h000;
            3555: color = 12'h000;
            3556: color = 12'h000;
            3557: color = 12'h000;
            3558: color = 12'h000;
            3559: color = 12'h000;
            3560: color = 12'h000;
            3561: color = 12'h000;
            3562: color = 12'h000;
            3563: color = 12'h000;
            3564: color = 12'h000;
            3565: color = 12'h000;
            3566: color = 12'h000;
            3567: color = 12'h000;
            3568: color = 12'h000;
            3569: color = 12'h000;
            3570: color = 12'h000;
            3571: color = 12'h000;
            3572: color = 12'h000;
            3573: color = 12'h000;
            3574: color = 12'h000;
            3575: color = 12'h000;
            3576: color = 12'h000;
            3577: color = 12'h000;
            3578: color = 12'h000;
            3579: color = 12'h000;
            3580: color = 12'h000;
            3581: color = 12'h000;
            3582: color = 12'h000;
            3583: color = 12'h000;
            3584: color = 12'h000;
            3585: color = 12'h000;
            3586: color = 12'h000;
            3587: color = 12'h000;
            3588: color = 12'h000;
            3589: color = 12'h000;
            3590: color = 12'h000;
            3591: color = 12'h000;
            3592: color = 12'h000;
            3593: color = 12'h000;
            3594: color = 12'h000;
            3595: color = 12'h000;
            3596: color = 12'h000;
            3597: color = 12'h000;
            3598: color = 12'h000;
            3599: color = 12'h000;
            3600: color = 12'h000;
            3601: color = 12'h000;
            3602: color = 12'h000;
            3603: color = 12'h000;
            3604: color = 12'h000;
            3605: color = 12'h000;
            3606: color = 12'h000;
            3607: color = 12'h000;
            3608: color = 12'h000;
            3609: color = 12'h000;
            3610: color = 12'h000;
            3611: color = 12'h000;
            3612: color = 12'h000;
            3613: color = 12'h000;
            3614: color = 12'h000;
            3615: color = 12'h000;
            3616: color = 12'h000;
            3617: color = 12'h000;
            3618: color = 12'h000;
            3619: color = 12'h000;
            3620: color = 12'h000;
            3621: color = 12'h000;
            3622: color = 12'h000;
            3623: color = 12'h000;
            3624: color = 12'h000;
            3625: color = 12'h000;
            3626: color = 12'h000;
            3627: color = 12'h000;
            3628: color = 12'h000;
            3629: color = 12'h000;
            3630: color = 12'h000;
            3631: color = 12'h000;
            3632: color = 12'h000;
            3633: color = 12'h000;
            3634: color = 12'h000;
            3635: color = 12'h000;
            3636: color = 12'h000;
            3637: color = 12'h000;
            3638: color = 12'h000;
            3639: color = 12'h000;
            3640: color = 12'h000;
            3641: color = 12'h000;
            3642: color = 12'h000;
            3643: color = 12'h000;
            3644: color = 12'h000;
            3645: color = 12'h000;
            3646: color = 12'h000;
            3647: color = 12'h000;
            3648: color = 12'h000;
            3649: color = 12'h000;
            3650: color = 12'h000;
            3651: color = 12'h000;
            3652: color = 12'h000;
            3653: color = 12'h000;
            3654: color = 12'h000;
            3655: color = 12'h000;
            3656: color = 12'h000;
            3657: color = 12'h000;
            3658: color = 12'h000;
            3659: color = 12'h000;
            3660: color = 12'h000;
            3661: color = 12'h000;
            3662: color = 12'h000;
            3663: color = 12'h000;
            3664: color = 12'h000;
            3665: color = 12'h000;
            3666: color = 12'h000;
            3667: color = 12'h000;
            3668: color = 12'h000;
            3669: color = 12'h000;
            3670: color = 12'h000;
            3671: color = 12'h000;
            3672: color = 12'h000;
            3673: color = 12'h000;
            3674: color = 12'h000;
            3675: color = 12'h000;
            3676: color = 12'h000;
            3677: color = 12'h000;
            3678: color = 12'h000;
            3679: color = 12'h000;
            3680: color = 12'h000;
            3681: color = 12'h000;
            3682: color = 12'h000;
            3683: color = 12'h000;
            3684: color = 12'h000;
            3685: color = 12'h000;
            3686: color = 12'h000;
            3687: color = 12'h000;
            3688: color = 12'h000;
            3689: color = 12'h000;
            3690: color = 12'h000;
            3691: color = 12'h000;
            3692: color = 12'h000;
            3693: color = 12'h000;
            3694: color = 12'h000;
            3695: color = 12'h000;
            3696: color = 12'h000;
            3697: color = 12'h000;
            3698: color = 12'h000;
            3699: color = 12'h000;
            3700: color = 12'h000;
            3701: color = 12'h000;
            3702: color = 12'h000;
            3703: color = 12'h000;
            3704: color = 12'h000;
            3705: color = 12'h000;
            3706: color = 12'h000;
            3707: color = 12'h000;
            3708: color = 12'h000;
            3709: color = 12'h000;
            3710: color = 12'h000;
            3711: color = 12'h000;
            3712: color = 12'h000;
            3713: color = 12'h000;
            3714: color = 12'h000;
            3715: color = 12'h000;
            3716: color = 12'h000;
            3717: color = 12'h000;
            3718: color = 12'h000;
            3719: color = 12'h000;
            3720: color = 12'h000;
            3721: color = 12'h000;
            3722: color = 12'h000;
            3723: color = 12'h000;
            3724: color = 12'h000;
            3725: color = 12'h000;
            3726: color = 12'h000;
            3727: color = 12'h000;
            3728: color = 12'h000;
            3729: color = 12'h000;
            3730: color = 12'h000;
            3731: color = 12'h000;
            3732: color = 12'h000;
            3733: color = 12'h000;
            3734: color = 12'h000;
            3735: color = 12'h000;
            3736: color = 12'h000;
            3737: color = 12'h000;
            3738: color = 12'h000;
            3739: color = 12'h000;
            3740: color = 12'h000;
            3741: color = 12'h000;
            3742: color = 12'h000;
            3743: color = 12'h000;
            3744: color = 12'h000;
            3745: color = 12'h000;
            3746: color = 12'h000;
            3747: color = 12'h000;
            3748: color = 12'h000;
            3749: color = 12'h000;
            3750: color = 12'h000;
            3751: color = 12'h000;
            3752: color = 12'h000;
            3753: color = 12'h000;
            3754: color = 12'h000;
            3755: color = 12'h000;
            3756: color = 12'h000;
            3757: color = 12'h000;
            3758: color = 12'h000;
            3759: color = 12'h000;
            3760: color = 12'h000;
            3761: color = 12'h000;
            3762: color = 12'h000;
            3763: color = 12'h000;
            3764: color = 12'h000;
            3765: color = 12'h000;
            3766: color = 12'h000;
            3767: color = 12'h000;
            3768: color = 12'h000;
            3769: color = 12'h000;
            3770: color = 12'h000;
            3771: color = 12'h000;
            3772: color = 12'h000;
            3773: color = 12'h000;
            3774: color = 12'h000;
            3775: color = 12'h000;
            3776: color = 12'h000;
            3777: color = 12'h000;
            3778: color = 12'h000;
            3779: color = 12'h000;
            3780: color = 12'h000;
            3781: color = 12'h000;
            3782: color = 12'h000;
            3783: color = 12'h000;
            3784: color = 12'h000;
            3785: color = 12'h000;
            3786: color = 12'h000;
            3787: color = 12'h000;
            3788: color = 12'h000;
            3789: color = 12'h000;
            3790: color = 12'h000;
            3791: color = 12'h000;
            3792: color = 12'h000;
            3793: color = 12'h000;
            3794: color = 12'h000;
            3795: color = 12'h000;
            3796: color = 12'h000;
            3797: color = 12'h000;
            3798: color = 12'h000;
            3799: color = 12'h000;
            3800: color = 12'h000;
            3801: color = 12'h000;
            3802: color = 12'h000;
            3803: color = 12'h000;
            3804: color = 12'h000;
            3805: color = 12'h000;
            3806: color = 12'h000;
            3807: color = 12'h000;
            3808: color = 12'h000;
            3809: color = 12'h000;
            3810: color = 12'h000;
            3811: color = 12'h000;
            3812: color = 12'h000;
            3813: color = 12'h000;
            3814: color = 12'h000;
            3815: color = 12'h000;
            3816: color = 12'h000;
            3817: color = 12'h000;
            3818: color = 12'h000;
            3819: color = 12'h000;
            3820: color = 12'h000;
            3821: color = 12'h000;
            3822: color = 12'h000;
            3823: color = 12'h000;
            3824: color = 12'h000;
            3825: color = 12'h000;
            3826: color = 12'h000;
            3827: color = 12'h000;
            3828: color = 12'h000;
            3829: color = 12'h000;
            3830: color = 12'h000;
            3831: color = 12'h000;
            3832: color = 12'h000;
            3833: color = 12'h000;
            3834: color = 12'h000;
            3835: color = 12'h000;
            3836: color = 12'h000;
            3837: color = 12'h000;
            3838: color = 12'h000;
            3839: color = 12'h000;
            3840: color = 12'h000;
            3841: color = 12'h000;
            3842: color = 12'h000;
            3843: color = 12'h000;
            3844: color = 12'h000;
            3845: color = 12'h000;
            3846: color = 12'h000;
            3847: color = 12'h000;
            3848: color = 12'h000;
            3849: color = 12'h000;
            3850: color = 12'h000;
            3851: color = 12'h000;
            3852: color = 12'h000;
            3853: color = 12'h000;
            3854: color = 12'h000;
            3855: color = 12'h000;
            3856: color = 12'h000;
            3857: color = 12'h000;
            3858: color = 12'h000;
            3859: color = 12'h000;
            3860: color = 12'h000;
            3861: color = 12'h000;
            3862: color = 12'h000;
            3863: color = 12'h000;
            3864: color = 12'h000;
            3865: color = 12'h000;
            3866: color = 12'h000;
            3867: color = 12'h000;
            3868: color = 12'h000;
            3869: color = 12'h000;
            3870: color = 12'h000;
            3871: color = 12'h000;
            3872: color = 12'h000;
            3873: color = 12'h000;
            3874: color = 12'h000;
            3875: color = 12'h000;
            3876: color = 12'h000;
            3877: color = 12'h000;
            3878: color = 12'h000;
            3879: color = 12'h000;
            3880: color = 12'h000;
            3881: color = 12'h000;
            3882: color = 12'h000;
            3883: color = 12'h000;
            3884: color = 12'h000;
            3885: color = 12'h000;
            3886: color = 12'h000;
            3887: color = 12'h000;
            3888: color = 12'h000;
            3889: color = 12'h000;
            3890: color = 12'h000;
            3891: color = 12'h000;
            3892: color = 12'h000;
            3893: color = 12'h000;
            3894: color = 12'h000;
            3895: color = 12'h000;
            3896: color = 12'h000;
            3897: color = 12'h000;
            3898: color = 12'h000;
            3899: color = 12'h000;
            3900: color = 12'h000;
            3901: color = 12'h000;
            3902: color = 12'h000;
            3903: color = 12'h000;
            3904: color = 12'h000;
            3905: color = 12'h000;
            3906: color = 12'h000;
            3907: color = 12'h000;
            3908: color = 12'h000;
            3909: color = 12'h000;
            3910: color = 12'h000;
            3911: color = 12'h000;
            3912: color = 12'h000;
            3913: color = 12'h000;
            3914: color = 12'h000;
            3915: color = 12'h000;
            3916: color = 12'h000;
            3917: color = 12'h000;
            3918: color = 12'h000;
            3919: color = 12'h000;
            3920: color = 12'h000;
            3921: color = 12'h000;
            3922: color = 12'h000;
            3923: color = 12'h000;
            3924: color = 12'h000;
            3925: color = 12'h000;
            3926: color = 12'h000;
            3927: color = 12'h000;
            3928: color = 12'h000;
            3929: color = 12'h000;
            3930: color = 12'h000;
            3931: color = 12'h000;
            3932: color = 12'h000;
            3933: color = 12'h000;
            3934: color = 12'h000;
            3935: color = 12'h000;
            3936: color = 12'h000;
            3937: color = 12'h000;
            3938: color = 12'h000;
            3939: color = 12'h000;
            3940: color = 12'h000;
            3941: color = 12'h000;
            3942: color = 12'h000;
            3943: color = 12'h000;
            3944: color = 12'h000;
            3945: color = 12'h000;
            3946: color = 12'h000;
            3947: color = 12'h000;
            3948: color = 12'h000;
            3949: color = 12'h000;
            3950: color = 12'h000;
            3951: color = 12'h000;
            3952: color = 12'h000;
            3953: color = 12'h000;
            3954: color = 12'h000;
            3955: color = 12'h000;
            3956: color = 12'h000;
            3957: color = 12'h000;
            3958: color = 12'h000;
            3959: color = 12'h000;
            3960: color = 12'h000;
            3961: color = 12'h000;
            3962: color = 12'h000;
            3963: color = 12'h000;
            3964: color = 12'h000;
            3965: color = 12'h000;
            3966: color = 12'h000;
            3967: color = 12'h000;
            3968: color = 12'h000;
            3969: color = 12'h000;
            3970: color = 12'h000;
            3971: color = 12'h000;
            3972: color = 12'h000;
            3973: color = 12'h000;
            3974: color = 12'h000;
            3975: color = 12'h000;
            3976: color = 12'h000;
            3977: color = 12'h000;
            3978: color = 12'h000;
            3979: color = 12'h000;
            3980: color = 12'h000;
            3981: color = 12'h000;
            3982: color = 12'h000;
            3983: color = 12'h000;
            3984: color = 12'h000;
            3985: color = 12'h000;
            3986: color = 12'h000;
            3987: color = 12'h000;
            3988: color = 12'h000;
            3989: color = 12'h000;
            3990: color = 12'h000;
            3991: color = 12'h000;
            3992: color = 12'h000;
            3993: color = 12'h000;
            3994: color = 12'h000;
            3995: color = 12'h000;
            3996: color = 12'h000;
            3997: color = 12'h000;
            3998: color = 12'h000;
            3999: color = 12'h000;
            4000: color = 12'h000;
            4001: color = 12'h000;
            4002: color = 12'h000;
            4003: color = 12'h000;
            4004: color = 12'h000;
            4005: color = 12'h000;
            4006: color = 12'h000;
            4007: color = 12'h000;
            4008: color = 12'h000;
            4009: color = 12'h000;
            4010: color = 12'h000;
            4011: color = 12'h000;
            4012: color = 12'h000;
            4013: color = 12'h000;
            4014: color = 12'h000;
            4015: color = 12'h000;
            4016: color = 12'h000;
            4017: color = 12'h000;
            4018: color = 12'h000;
            4019: color = 12'h000;
            4020: color = 12'h000;
            4021: color = 12'h000;
            4022: color = 12'h000;
            4023: color = 12'h000;
            4024: color = 12'h000;
            4025: color = 12'h000;
            4026: color = 12'h000;
            4027: color = 12'h000;
            4028: color = 12'h000;
            4029: color = 12'h000;
            4030: color = 12'h000;
            4031: color = 12'h000;
            4032: color = 12'h000;
            4033: color = 12'h000;
            4034: color = 12'h000;
            4035: color = 12'h000;
            4036: color = 12'h000;
            4037: color = 12'h000;
            4038: color = 12'h000;
            4039: color = 12'h000;
            4040: color = 12'h000;
            4041: color = 12'h000;
            4042: color = 12'h000;
            4043: color = 12'h000;
            4044: color = 12'h000;
            4045: color = 12'h000;
            4046: color = 12'h000;
            4047: color = 12'h000;
            4048: color = 12'h000;
            4049: color = 12'h000;
            4050: color = 12'h000;
            4051: color = 12'h000;
            4052: color = 12'h000;
            4053: color = 12'h000;
            4054: color = 12'h000;
            4055: color = 12'h000;
            4056: color = 12'h000;
            4057: color = 12'h000;
            4058: color = 12'h000;
            4059: color = 12'h000;
            4060: color = 12'h000;
            4061: color = 12'h000;
            4062: color = 12'h000;
            4063: color = 12'h000;
            4064: color = 12'h000;
            4065: color = 12'h000;
            4066: color = 12'h000;
            4067: color = 12'h000;
            4068: color = 12'h000;
            4069: color = 12'h000;
            4070: color = 12'h000;
            4071: color = 12'h000;
            4072: color = 12'h000;
            4073: color = 12'h000;
            4074: color = 12'h000;
            4075: color = 12'h000;
            4076: color = 12'h000;
            4077: color = 12'h000;
            4078: color = 12'h000;
            4079: color = 12'h000;
            4080: color = 12'h000;
            4081: color = 12'h000;
            4082: color = 12'h000;
            4083: color = 12'h000;
            4084: color = 12'h000;
            4085: color = 12'h000;
            4086: color = 12'h000;
            4087: color = 12'h000;
            4088: color = 12'h000;
            4089: color = 12'h000;
            4090: color = 12'h000;
            4091: color = 12'h000;
            4092: color = 12'h000;
            4093: color = 12'h000;
            4094: color = 12'h000;
            4095: color = 12'h000;
            4096: color = 12'h000;
            4097: color = 12'h000;
            4098: color = 12'h000;
            4099: color = 12'h000;
            4100: color = 12'h000;
            4101: color = 12'h000;
            4102: color = 12'h000;
            4103: color = 12'h000;
            4104: color = 12'h000;
            4105: color = 12'h000;
            4106: color = 12'h000;
            4107: color = 12'h000;
            4108: color = 12'h000;
            4109: color = 12'h000;
            4110: color = 12'h000;
            4111: color = 12'h000;
            4112: color = 12'h000;
            4113: color = 12'h000;
            4114: color = 12'h000;
            4115: color = 12'h000;
            4116: color = 12'h000;
            4117: color = 12'h000;
            4118: color = 12'h000;
            4119: color = 12'h000;
            4120: color = 12'h000;
            4121: color = 12'h000;
            4122: color = 12'h000;
            4123: color = 12'h000;
            4124: color = 12'h000;
            4125: color = 12'h000;
            4126: color = 12'h000;
            4127: color = 12'h000;
            4128: color = 12'h000;
            4129: color = 12'h000;
            4130: color = 12'h000;
            4131: color = 12'h000;
            4132: color = 12'h000;
            4133: color = 12'h000;
            4134: color = 12'h000;
            4135: color = 12'h000;
            4136: color = 12'h000;
            4137: color = 12'h000;
            4138: color = 12'h000;
            4139: color = 12'h000;
            4140: color = 12'h000;
            4141: color = 12'h000;
            4142: color = 12'h000;
            4143: color = 12'h000;
            4144: color = 12'h000;
            4145: color = 12'h000;
            4146: color = 12'h000;
            4147: color = 12'h000;
            4148: color = 12'h000;
            4149: color = 12'h000;
            4150: color = 12'h000;
            4151: color = 12'h000;
            4152: color = 12'h000;
            4153: color = 12'h000;
            4154: color = 12'h000;
            4155: color = 12'h000;
            4156: color = 12'h000;
            4157: color = 12'h000;
            4158: color = 12'h000;
            4159: color = 12'h000;
            4160: color = 12'h000;
            4161: color = 12'h000;
            4162: color = 12'h000;
            4163: color = 12'h000;
            4164: color = 12'h000;
            4165: color = 12'h000;
            4166: color = 12'h000;
            4167: color = 12'h000;
            4168: color = 12'h000;
            4169: color = 12'h000;
            4170: color = 12'h000;
            4171: color = 12'h000;
            4172: color = 12'h000;
            4173: color = 12'h000;
            4174: color = 12'h000;
            4175: color = 12'h000;
            4176: color = 12'h000;
            4177: color = 12'h000;
            4178: color = 12'h000;
            4179: color = 12'h000;
            4180: color = 12'h000;
            4181: color = 12'h000;
            4182: color = 12'h000;
            4183: color = 12'h000;
            4184: color = 12'h000;
            4185: color = 12'h000;
            4186: color = 12'h000;
            4187: color = 12'h000;
            4188: color = 12'h000;
            4189: color = 12'h000;
            4190: color = 12'h000;
            4191: color = 12'h000;
            4192: color = 12'h000;
            4193: color = 12'h000;
            4194: color = 12'h000;
            4195: color = 12'h000;
            4196: color = 12'h000;
            4197: color = 12'h000;
            4198: color = 12'h000;
            4199: color = 12'h000;
            4200: color = 12'h000;
            4201: color = 12'h000;
            4202: color = 12'h000;
            4203: color = 12'h000;
            4204: color = 12'h000;
            4205: color = 12'h000;
            4206: color = 12'h000;
            4207: color = 12'h000;
            4208: color = 12'h000;
            4209: color = 12'h000;
            4210: color = 12'h000;
            4211: color = 12'h000;
            4212: color = 12'h000;
            4213: color = 12'h000;
            4214: color = 12'h000;
            4215: color = 12'h000;
            4216: color = 12'h000;
            4217: color = 12'h000;
            4218: color = 12'h000;
            4219: color = 12'h000;
            4220: color = 12'h000;
            4221: color = 12'h000;
            4222: color = 12'h000;
            4223: color = 12'h000;
            4224: color = 12'h000;
            4225: color = 12'h000;
            4226: color = 12'h000;
            4227: color = 12'h000;
            4228: color = 12'h000;
            4229: color = 12'h000;
            4230: color = 12'h000;
            4231: color = 12'h000;
            4232: color = 12'h000;
            4233: color = 12'h000;
            4234: color = 12'h000;
            4235: color = 12'h000;
            4236: color = 12'h000;
            4237: color = 12'h000;
            4238: color = 12'h000;
            4239: color = 12'h000;
            4240: color = 12'h000;
            4241: color = 12'h000;
            4242: color = 12'h000;
            4243: color = 12'h000;
            4244: color = 12'h000;
            4245: color = 12'h000;
            4246: color = 12'h000;
            4247: color = 12'h000;
            4248: color = 12'h000;
            4249: color = 12'h000;
            4250: color = 12'h000;
            4251: color = 12'h000;
            4252: color = 12'h000;
            4253: color = 12'h000;
            4254: color = 12'h000;
            4255: color = 12'h000;
            4256: color = 12'h000;
            4257: color = 12'h000;
            4258: color = 12'h000;
            4259: color = 12'h000;
            4260: color = 12'h000;
            4261: color = 12'h000;
            4262: color = 12'h000;
            4263: color = 12'h000;
            4264: color = 12'h000;
            4265: color = 12'h000;
            4266: color = 12'h000;
            4267: color = 12'h000;
            4268: color = 12'h000;
            4269: color = 12'h000;
            4270: color = 12'h000;
            4271: color = 12'h000;
            4272: color = 12'h000;
            4273: color = 12'h000;
            4274: color = 12'h000;
            4275: color = 12'h000;
            4276: color = 12'h000;
            4277: color = 12'h000;
            4278: color = 12'h000;
            4279: color = 12'h000;
            4280: color = 12'h000;
            4281: color = 12'h000;
            4282: color = 12'h000;
            4283: color = 12'h000;
            4284: color = 12'h000;
            4285: color = 12'h000;
            4286: color = 12'h000;
            4287: color = 12'h000;
            4288: color = 12'h000;
            4289: color = 12'h000;
            4290: color = 12'h000;
            4291: color = 12'h000;
            4292: color = 12'h000;
            4293: color = 12'h000;
            4294: color = 12'h000;
            4295: color = 12'h000;
            4296: color = 12'h000;
            4297: color = 12'h000;
            4298: color = 12'h000;
            4299: color = 12'h000;
            4300: color = 12'h000;
            4301: color = 12'h000;
            4302: color = 12'h000;
            4303: color = 12'h000;
            4304: color = 12'h000;
            4305: color = 12'h000;
            4306: color = 12'h000;
            4307: color = 12'h000;
            4308: color = 12'h000;
            4309: color = 12'h000;
            4310: color = 12'h000;
            4311: color = 12'h000;
            4312: color = 12'h000;
            4313: color = 12'h000;
            4314: color = 12'h000;
            4315: color = 12'h000;
            4316: color = 12'h000;
            4317: color = 12'h000;
            4318: color = 12'h000;
            4319: color = 12'h000;
            4320: color = 12'h000;
            4321: color = 12'h000;
            4322: color = 12'h000;
            4323: color = 12'h000;
            4324: color = 12'h000;
            4325: color = 12'h000;
            4326: color = 12'h000;
            4327: color = 12'h000;
            4328: color = 12'h000;
            4329: color = 12'h000;
            4330: color = 12'h000;
            4331: color = 12'h000;
            4332: color = 12'h000;
            4333: color = 12'h000;
            4334: color = 12'h000;
            4335: color = 12'h000;
            4336: color = 12'h000;
            4337: color = 12'h000;
            4338: color = 12'h000;
            4339: color = 12'h000;
            4340: color = 12'h000;
            4341: color = 12'h000;
            4342: color = 12'h000;
            4343: color = 12'h000;
            4344: color = 12'h000;
            4345: color = 12'h000;
            4346: color = 12'h000;
            4347: color = 12'h000;
            4348: color = 12'h000;
            4349: color = 12'h000;
            4350: color = 12'h000;
            4351: color = 12'h000;
            4352: color = 12'h000;
            4353: color = 12'h000;
            4354: color = 12'h000;
            4355: color = 12'h000;
            4356: color = 12'h000;
            4357: color = 12'h000;
            4358: color = 12'h000;
            4359: color = 12'h000;
            4360: color = 12'h000;
            4361: color = 12'h000;
            4362: color = 12'h000;
            4363: color = 12'h000;
            4364: color = 12'h000;
            4365: color = 12'h000;
            4366: color = 12'h000;
            4367: color = 12'h000;
            4368: color = 12'h000;
            4369: color = 12'h000;
            4370: color = 12'h000;
            4371: color = 12'h000;
            4372: color = 12'h000;
            4373: color = 12'h000;
            4374: color = 12'h000;
            4375: color = 12'h000;
            4376: color = 12'h000;
            4377: color = 12'h000;
            4378: color = 12'h000;
            4379: color = 12'h000;
            4380: color = 12'h000;
            4381: color = 12'h000;
            4382: color = 12'h000;
            4383: color = 12'h000;
            4384: color = 12'h000;
            4385: color = 12'h000;
            4386: color = 12'h000;
            4387: color = 12'h000;
            4388: color = 12'h000;
            4389: color = 12'h000;
            4390: color = 12'h000;
            4391: color = 12'h000;
            4392: color = 12'h000;
            4393: color = 12'h000;
            4394: color = 12'h000;
            4395: color = 12'h000;
            4396: color = 12'h000;
            4397: color = 12'h000;
            4398: color = 12'h000;
            4399: color = 12'h000;
            4400: color = 12'h000;
            4401: color = 12'h000;
            4402: color = 12'h000;
            4403: color = 12'h000;
            4404: color = 12'h000;
            4405: color = 12'h000;
            4406: color = 12'h000;
            4407: color = 12'h000;
            4408: color = 12'h000;
            4409: color = 12'h000;
            4410: color = 12'h000;
            4411: color = 12'h000;
            4412: color = 12'h000;
            4413: color = 12'h000;
            4414: color = 12'h000;
            4415: color = 12'h000;
            4416: color = 12'h000;
            4417: color = 12'h000;
            4418: color = 12'h000;
            4419: color = 12'h000;
            4420: color = 12'h000;
            4421: color = 12'h000;
            4422: color = 12'h000;
            4423: color = 12'h000;
            4424: color = 12'h000;
            4425: color = 12'h000;
            4426: color = 12'h000;
            4427: color = 12'h000;
            4428: color = 12'h000;
            4429: color = 12'h000;
            4430: color = 12'h000;
            4431: color = 12'h000;
            4432: color = 12'h000;
            4433: color = 12'h000;
            4434: color = 12'h000;
            4435: color = 12'h000;
            4436: color = 12'h000;
            4437: color = 12'h000;
            4438: color = 12'h000;
            4439: color = 12'h000;
            4440: color = 12'h000;
            4441: color = 12'h000;
            4442: color = 12'h000;
            4443: color = 12'h000;
            4444: color = 12'h000;
            4445: color = 12'h000;
            4446: color = 12'h000;
            4447: color = 12'h000;
            4448: color = 12'h000;
            4449: color = 12'h000;
            4450: color = 12'h000;
            4451: color = 12'h000;
            4452: color = 12'h000;
            4453: color = 12'h000;
            4454: color = 12'h000;
            4455: color = 12'h000;
            4456: color = 12'h000;
            4457: color = 12'h000;
            4458: color = 12'h000;
            4459: color = 12'h000;
            4460: color = 12'h000;
            4461: color = 12'h000;
            4462: color = 12'h000;
            4463: color = 12'h000;
            4464: color = 12'h000;
            4465: color = 12'h000;
            4466: color = 12'h000;
            4467: color = 12'h000;
            4468: color = 12'h000;
            4469: color = 12'h000;
            4470: color = 12'h000;
            4471: color = 12'h000;
            4472: color = 12'h000;
            4473: color = 12'h000;
            4474: color = 12'h000;
            4475: color = 12'h000;
            4476: color = 12'h000;
            4477: color = 12'h000;
            4478: color = 12'h000;
            4479: color = 12'h000;
            4480: color = 12'h000;
            4481: color = 12'h000;
            4482: color = 12'h000;
            4483: color = 12'h000;
            4484: color = 12'h000;
            4485: color = 12'h000;
            4486: color = 12'h000;
            4487: color = 12'h000;
            4488: color = 12'h000;
            4489: color = 12'h000;
            4490: color = 12'h000;
            4491: color = 12'h000;
            4492: color = 12'h000;
            4493: color = 12'h000;
            4494: color = 12'h000;
            4495: color = 12'h000;
            4496: color = 12'h000;
            4497: color = 12'h000;
            4498: color = 12'h000;
            4499: color = 12'h000;
            4500: color = 12'h000;
            4501: color = 12'h000;
            4502: color = 12'h000;
            4503: color = 12'h000;
            4504: color = 12'h000;
            4505: color = 12'h000;
            4506: color = 12'h000;
            4507: color = 12'h000;
            4508: color = 12'h000;
            4509: color = 12'h000;
            4510: color = 12'h000;
            4511: color = 12'h000;
            4512: color = 12'h000;
            4513: color = 12'h000;
            4514: color = 12'h000;
            4515: color = 12'h000;
            4516: color = 12'h000;
            4517: color = 12'h000;
            4518: color = 12'h000;
            4519: color = 12'h000;
            4520: color = 12'h000;
            4521: color = 12'h000;
            4522: color = 12'h000;
            4523: color = 12'h000;
            4524: color = 12'h000;
            4525: color = 12'h000;
            4526: color = 12'h000;
            4527: color = 12'h000;
            4528: color = 12'h000;
            4529: color = 12'h000;
            4530: color = 12'h000;
            4531: color = 12'h000;
            4532: color = 12'h000;
            4533: color = 12'h000;
            4534: color = 12'h000;
            4535: color = 12'h000;
            4536: color = 12'h000;
            4537: color = 12'h000;
            4538: color = 12'h000;
            4539: color = 12'h000;
            4540: color = 12'h000;
            4541: color = 12'h000;
            4542: color = 12'h000;
            4543: color = 12'h000;
            4544: color = 12'h000;
            4545: color = 12'h000;
            4546: color = 12'h000;
            4547: color = 12'h000;
            4548: color = 12'h000;
            4549: color = 12'h000;
            4550: color = 12'h000;
            4551: color = 12'h000;
            4552: color = 12'h000;
            4553: color = 12'h000;
            4554: color = 12'h000;
            4555: color = 12'h000;
            4556: color = 12'h000;
            4557: color = 12'h000;
            4558: color = 12'h000;
            4559: color = 12'h000;
            4560: color = 12'h000;
            4561: color = 12'h000;
            4562: color = 12'h000;
            4563: color = 12'h000;
            4564: color = 12'h000;
            4565: color = 12'h000;
            4566: color = 12'h000;
            4567: color = 12'h000;
            4568: color = 12'h000;
            4569: color = 12'h000;
            4570: color = 12'h000;
            4571: color = 12'h000;
            4572: color = 12'h000;
            4573: color = 12'h000;
            4574: color = 12'h000;
            4575: color = 12'h000;
            4576: color = 12'h000;
            4577: color = 12'h000;
            4578: color = 12'h000;
            4579: color = 12'h000;
            4580: color = 12'h000;
            4581: color = 12'h000;
            4582: color = 12'h000;
            4583: color = 12'h000;
            4584: color = 12'h000;
            4585: color = 12'h000;
            4586: color = 12'h000;
            4587: color = 12'h000;
            4588: color = 12'h000;
            4589: color = 12'h000;
            4590: color = 12'h000;
            4591: color = 12'h000;
            4592: color = 12'h000;
            4593: color = 12'h000;
            4594: color = 12'h000;
            4595: color = 12'h000;
            4596: color = 12'h000;
            4597: color = 12'h000;
            4598: color = 12'h000;
            4599: color = 12'h000;
            4600: color = 12'h000;
            4601: color = 12'h000;
            4602: color = 12'h000;
            4603: color = 12'h000;
            4604: color = 12'h000;
            4605: color = 12'h000;
            4606: color = 12'h000;
            4607: color = 12'h000;
            4608: color = 12'h000;
            4609: color = 12'h000;
            4610: color = 12'h000;
            4611: color = 12'h000;
            4612: color = 12'h000;
            4613: color = 12'h000;
            4614: color = 12'h000;
            4615: color = 12'h000;
            4616: color = 12'h000;
            4617: color = 12'h000;
            4618: color = 12'h000;
            4619: color = 12'h000;
            4620: color = 12'h000;
            4621: color = 12'h000;
            4622: color = 12'h000;
            4623: color = 12'h000;
            4624: color = 12'h000;
            4625: color = 12'h000;
            4626: color = 12'h000;
            4627: color = 12'h000;
            4628: color = 12'h000;
            4629: color = 12'h000;
            4630: color = 12'h000;
            4631: color = 12'h000;
            4632: color = 12'h000;
            4633: color = 12'h000;
            4634: color = 12'h000;
            4635: color = 12'h000;
            4636: color = 12'h000;
            4637: color = 12'h000;
            4638: color = 12'h000;
            4639: color = 12'h000;
            4640: color = 12'h000;
            4641: color = 12'h000;
            4642: color = 12'h000;
            4643: color = 12'h000;
            4644: color = 12'h000;
            4645: color = 12'h000;
            4646: color = 12'h000;
            4647: color = 12'h000;
            4648: color = 12'h000;
            4649: color = 12'h000;
            4650: color = 12'h000;
            4651: color = 12'h000;
            4652: color = 12'h000;
            4653: color = 12'h000;
            4654: color = 12'h000;
            4655: color = 12'h000;
            4656: color = 12'h000;
            4657: color = 12'h000;
            4658: color = 12'h000;
            4659: color = 12'h000;
            4660: color = 12'h000;
            4661: color = 12'h000;
            4662: color = 12'h000;
            4663: color = 12'h000;
            4664: color = 12'h000;
            4665: color = 12'h000;
            4666: color = 12'h000;
            4667: color = 12'h000;
            4668: color = 12'h000;
            4669: color = 12'h000;
            4670: color = 12'h000;
            4671: color = 12'h000;
            4672: color = 12'h000;
            4673: color = 12'h000;
            4674: color = 12'h000;
            4675: color = 12'h000;
            4676: color = 12'h000;
            4677: color = 12'h000;
            4678: color = 12'h000;
            4679: color = 12'h000;
            4680: color = 12'h000;
            4681: color = 12'h000;
            4682: color = 12'h000;
            4683: color = 12'h000;
            4684: color = 12'h000;
            4685: color = 12'h000;
            4686: color = 12'h000;
            4687: color = 12'h000;
            4688: color = 12'h000;
            4689: color = 12'h000;
            4690: color = 12'h000;
            4691: color = 12'h000;
            4692: color = 12'h000;
            4693: color = 12'h000;
            4694: color = 12'h000;
            4695: color = 12'h000;
            4696: color = 12'h000;
            4697: color = 12'h000;
            4698: color = 12'h000;
            4699: color = 12'h000;
            4700: color = 12'h000;
            4701: color = 12'h000;
            4702: color = 12'h000;
            4703: color = 12'h000;
            4704: color = 12'h000;
            4705: color = 12'h000;
            4706: color = 12'h000;
            4707: color = 12'h000;
            4708: color = 12'h000;
            4709: color = 12'h000;
            4710: color = 12'h000;
            4711: color = 12'h000;
            4712: color = 12'h000;
            4713: color = 12'h000;
            4714: color = 12'h000;
            4715: color = 12'h000;
            4716: color = 12'h000;
            4717: color = 12'h000;
            4718: color = 12'h000;
            4719: color = 12'h000;
            4720: color = 12'h000;
            4721: color = 12'h000;
            4722: color = 12'h000;
            4723: color = 12'h000;
            4724: color = 12'h000;
            4725: color = 12'h000;
            4726: color = 12'h000;
            4727: color = 12'h000;
            4728: color = 12'h000;
            4729: color = 12'h000;
            4730: color = 12'h000;
            4731: color = 12'h000;
            4732: color = 12'h000;
            4733: color = 12'h000;
            4734: color = 12'h000;
            4735: color = 12'h000;
            4736: color = 12'h000;
            4737: color = 12'h000;
            4738: color = 12'h000;
            4739: color = 12'h000;
            4740: color = 12'h000;
            4741: color = 12'h000;
            4742: color = 12'h000;
            4743: color = 12'h000;
            4744: color = 12'h000;
            4745: color = 12'h000;
            4746: color = 12'h000;
            4747: color = 12'h000;
            4748: color = 12'h000;
            4749: color = 12'h000;
            4750: color = 12'h000;
            4751: color = 12'h000;
            4752: color = 12'h000;
            4753: color = 12'h000;
            4754: color = 12'h000;
            4755: color = 12'h000;
            4756: color = 12'h000;
            4757: color = 12'h000;
            4758: color = 12'h000;
            4759: color = 12'h000;
            4760: color = 12'h000;
            4761: color = 12'h000;
            4762: color = 12'h000;
            4763: color = 12'h000;
            4764: color = 12'h000;
            4765: color = 12'h000;
            4766: color = 12'h000;
            4767: color = 12'h000;
            4768: color = 12'h000;
            4769: color = 12'h000;
            4770: color = 12'h000;
            4771: color = 12'h000;
            4772: color = 12'h000;
            4773: color = 12'h000;
            4774: color = 12'h000;
            4775: color = 12'h000;
            4776: color = 12'h000;
            4777: color = 12'h000;
            4778: color = 12'h000;
            4779: color = 12'h000;
            4780: color = 12'h000;
            4781: color = 12'h000;
            4782: color = 12'h000;
            4783: color = 12'h000;
            4784: color = 12'h000;
            4785: color = 12'h000;
            4786: color = 12'h000;
            4787: color = 12'h000;
            4788: color = 12'h000;
            4789: color = 12'h000;
            4790: color = 12'h000;
            4791: color = 12'h000;
            4792: color = 12'h000;
            4793: color = 12'h000;
            4794: color = 12'h000;
            4795: color = 12'h000;
            4796: color = 12'h000;
            4797: color = 12'h000;
            4798: color = 12'h000;
            4799: color = 12'h000;
            4800: color = 12'h000;
            4801: color = 12'h000;
            4802: color = 12'h000;
            4803: color = 12'h000;
            4804: color = 12'h000;
            4805: color = 12'h000;
            4806: color = 12'h000;
            4807: color = 12'h000;
            4808: color = 12'h000;
            4809: color = 12'h000;
            4810: color = 12'h000;
            4811: color = 12'h000;
            4812: color = 12'h000;
            4813: color = 12'h000;
            4814: color = 12'h000;
            4815: color = 12'h000;
            4816: color = 12'h000;
            4817: color = 12'h000;
            4818: color = 12'h000;
            4819: color = 12'h000;
            4820: color = 12'h000;
            4821: color = 12'h000;
            4822: color = 12'h000;
            4823: color = 12'h000;
            4824: color = 12'h000;
            4825: color = 12'h000;
            4826: color = 12'h000;
            4827: color = 12'h000;
            4828: color = 12'h000;
            4829: color = 12'h000;
            4830: color = 12'h000;
            4831: color = 12'h000;
            4832: color = 12'h000;
            4833: color = 12'h000;
            4834: color = 12'h000;
            4835: color = 12'h000;
            4836: color = 12'h000;
            4837: color = 12'h000;
            4838: color = 12'h000;
            4839: color = 12'h000;
            4840: color = 12'h000;
            4841: color = 12'h000;
            4842: color = 12'h000;
            4843: color = 12'h000;
            4844: color = 12'h000;
            4845: color = 12'h000;
            4846: color = 12'h000;
            4847: color = 12'h000;
            4848: color = 12'h000;
            4849: color = 12'h777;
            4850: color = 12'hFFF;
            4851: color = 12'hFFF;
            4852: color = 12'hFFF;
            4853: color = 12'hFFF;
            4854: color = 12'hFFF;
            4855: color = 12'hFFF;
            4856: color = 12'hFFF;
            4857: color = 12'hFFF;
            4858: color = 12'hFFF;
            4859: color = 12'hFFF;
            4860: color = 12'hFFF;
            4861: color = 12'h777;
            4862: color = 12'h000;
            4863: color = 12'h000;
            4864: color = 12'h000;
            4865: color = 12'h000;
            4866: color = 12'h000;
            4867: color = 12'h000;
            4868: color = 12'h000;
            4869: color = 12'h000;
            4870: color = 12'h000;
            4871: color = 12'h000;
            4872: color = 12'h000;
            4873: color = 12'h000;
            4874: color = 12'h000;
            4875: color = 12'h000;
            4876: color = 12'h000;
            4877: color = 12'h000;
            4878: color = 12'h000;
            4879: color = 12'h000;
            4880: color = 12'h000;
            4881: color = 12'h000;
            4882: color = 12'h000;
            4883: color = 12'h000;
            4884: color = 12'h000;
            4885: color = 12'h000;
            4886: color = 12'h000;
            4887: color = 12'h000;
            4888: color = 12'h000;
            4889: color = 12'h000;
            4890: color = 12'h000;
            4891: color = 12'h000;
            4892: color = 12'h000;
            4893: color = 12'h000;
            4894: color = 12'h000;
            4895: color = 12'h000;
            4896: color = 12'h000;
            4897: color = 12'h000;
            4898: color = 12'h000;
            4899: color = 12'h000;
            4900: color = 12'h000;
            4901: color = 12'h000;
            4902: color = 12'h000;
            4903: color = 12'h000;
            4904: color = 12'h000;
            4905: color = 12'h000;
            4906: color = 12'h000;
            4907: color = 12'h000;
            4908: color = 12'h000;
            4909: color = 12'h000;
            4910: color = 12'h000;
            4911: color = 12'h000;
            4912: color = 12'h000;
            4913: color = 12'h000;
            4914: color = 12'h000;
            4915: color = 12'h000;
            4916: color = 12'h000;
            4917: color = 12'h000;
            4918: color = 12'h000;
            4919: color = 12'h000;
            4920: color = 12'h000;
            4921: color = 12'h000;
            4922: color = 12'h000;
            4923: color = 12'hEEE;
            4924: color = 12'hFFF;
            4925: color = 12'hFFF;
            4926: color = 12'hFFF;
            4927: color = 12'hFFF;
            4928: color = 12'hFFF;
            4929: color = 12'hFFF;
            4930: color = 12'hFFF;
            4931: color = 12'hFFF;
            4932: color = 12'hFFF;
            4933: color = 12'hFFF;
            4934: color = 12'hFFF;
            4935: color = 12'hFFF;
            4936: color = 12'hFFF;
            4937: color = 12'hEEE;
            4938: color = 12'h000;
            4939: color = 12'h000;
            4940: color = 12'h000;
            4941: color = 12'h000;
            4942: color = 12'h000;
            4943: color = 12'h000;
            4944: color = 12'h000;
            4945: color = 12'h000;
            4946: color = 12'h000;
            4947: color = 12'h000;
            4948: color = 12'h000;
            4949: color = 12'h000;
            4950: color = 12'h000;
            4951: color = 12'h000;
            4952: color = 12'h000;
            4953: color = 12'h000;
            4954: color = 12'h000;
            4955: color = 12'h000;
            4956: color = 12'h000;
            4957: color = 12'h000;
            4958: color = 12'h000;
            4959: color = 12'h000;
            4960: color = 12'h000;
            4961: color = 12'h000;
            4962: color = 12'h000;
            4963: color = 12'h000;
            4964: color = 12'h000;
            4965: color = 12'h000;
            4966: color = 12'h000;
            4967: color = 12'h000;
            4968: color = 12'h000;
            4969: color = 12'h000;
            4970: color = 12'h000;
            4971: color = 12'h000;
            4972: color = 12'h000;
            4973: color = 12'h000;
            4974: color = 12'h000;
            4975: color = 12'h000;
            4976: color = 12'h000;
            4977: color = 12'h000;
            4978: color = 12'h000;
            4979: color = 12'h000;
            4980: color = 12'h000;
            4981: color = 12'h000;
            4982: color = 12'h000;
            4983: color = 12'h000;
            4984: color = 12'h000;
            4985: color = 12'h000;
            4986: color = 12'h000;
            4987: color = 12'h000;
            4988: color = 12'h000;
            4989: color = 12'h000;
            4990: color = 12'h000;
            4991: color = 12'h000;
            4992: color = 12'h000;
            4993: color = 12'h000;
            4994: color = 12'h000;
            4995: color = 12'h000;
            4996: color = 12'h000;
            4997: color = 12'h000;
            4998: color = 12'h000;
            4999: color = 12'h000;
            5000: color = 12'h000;
            5001: color = 12'h000;
            5002: color = 12'h000;
            5003: color = 12'h000;
            5004: color = 12'h000;
            5005: color = 12'h000;
            5006: color = 12'h000;
            5007: color = 12'h000;
            5008: color = 12'h000;
            5009: color = 12'h000;
            5010: color = 12'h000;
            5011: color = 12'h000;
            5012: color = 12'h000;
            5013: color = 12'h000;
            5014: color = 12'h000;
            5015: color = 12'h000;
            5016: color = 12'h000;
            5017: color = 12'h000;
            5018: color = 12'h000;
            5019: color = 12'h000;
            5020: color = 12'h000;
            5021: color = 12'h000;
            5022: color = 12'h000;
            5023: color = 12'h000;
            5024: color = 12'h000;
            5025: color = 12'h000;
            5026: color = 12'h000;
            5027: color = 12'h000;
            5028: color = 12'h000;
            5029: color = 12'h777;
            5030: color = 12'hFFF;
            5031: color = 12'hFFF;
            5032: color = 12'hFFF;
            5033: color = 12'hFFF;
            5034: color = 12'hFFF;
            5035: color = 12'hFFF;
            5036: color = 12'hFFF;
            5037: color = 12'hFFF;
            5038: color = 12'hFFF;
            5039: color = 12'hEEE;
            5040: color = 12'h000;
            5041: color = 12'h000;
            5042: color = 12'h000;
            5043: color = 12'h000;
            5044: color = 12'h000;
            5045: color = 12'h000;
            5046: color = 12'h000;
            5047: color = 12'h000;
            5048: color = 12'h000;
            5049: color = 12'h000;
            5050: color = 12'h000;
            5051: color = 12'h000;
            5052: color = 12'h000;
            5053: color = 12'h000;
            5054: color = 12'h000;
            5055: color = 12'h000;
            5056: color = 12'h000;
            5057: color = 12'h000;
            5058: color = 12'h000;
            5059: color = 12'h000;
            5060: color = 12'h000;
            5061: color = 12'h000;
            5062: color = 12'h000;
            5063: color = 12'h000;
            5064: color = 12'h000;
            5065: color = 12'h000;
            5066: color = 12'h000;
            5067: color = 12'h000;
            5068: color = 12'h000;
            5069: color = 12'h000;
            5070: color = 12'h000;
            5071: color = 12'h000;
            5072: color = 12'h000;
            5073: color = 12'h000;
            5074: color = 12'h000;
            5075: color = 12'h000;
            5076: color = 12'h000;
            5077: color = 12'h000;
            5078: color = 12'h000;
            5079: color = 12'h000;
            5080: color = 12'h000;
            5081: color = 12'h000;
            5082: color = 12'h000;
            5083: color = 12'h000;
            5084: color = 12'h000;
            5085: color = 12'h000;
            5086: color = 12'h000;
            5087: color = 12'h000;
            5088: color = 12'h000;
            5089: color = 12'h000;
            5090: color = 12'h000;
            5091: color = 12'h000;
            5092: color = 12'h000;
            5093: color = 12'h000;
            5094: color = 12'h000;
            5095: color = 12'h000;
            5096: color = 12'h000;
            5097: color = 12'h000;
            5098: color = 12'h000;
            5099: color = 12'h000;
            5100: color = 12'h000;
            5101: color = 12'h000;
            5102: color = 12'h000;
            5103: color = 12'h000;
            5104: color = 12'h000;
            5105: color = 12'h000;
            5106: color = 12'h000;
            5107: color = 12'h000;
            5108: color = 12'h000;
            5109: color = 12'h000;
            5110: color = 12'h000;
            5111: color = 12'h000;
            5112: color = 12'h000;
            5113: color = 12'h000;
            5114: color = 12'h000;
            5115: color = 12'h000;
            5116: color = 12'h000;
            5117: color = 12'h000;
            5118: color = 12'h000;
            5119: color = 12'h000;
            5120: color = 12'h000;
            5121: color = 12'h000;
            5122: color = 12'h000;
            5123: color = 12'h000;
            5124: color = 12'h000;
            5125: color = 12'h000;
            5126: color = 12'h000;
            5127: color = 12'h000;
            5128: color = 12'h000;
            5129: color = 12'h000;
            5130: color = 12'h000;
            5131: color = 12'h000;
            5132: color = 12'h000;
            5133: color = 12'h000;
            5134: color = 12'h000;
            5135: color = 12'h000;
            5136: color = 12'h000;
            5137: color = 12'h000;
            5138: color = 12'h000;
            5139: color = 12'h000;
            5140: color = 12'h000;
            5141: color = 12'h000;
            5142: color = 12'h000;
            5143: color = 12'h000;
            5144: color = 12'h000;
            5145: color = 12'h000;
            5146: color = 12'h000;
            5147: color = 12'h000;
            5148: color = 12'h000;
            5149: color = 12'h000;
            5150: color = 12'h000;
            5151: color = 12'h000;
            5152: color = 12'h000;
            5153: color = 12'h000;
            5154: color = 12'h000;
            5155: color = 12'h000;
            5156: color = 12'h000;
            5157: color = 12'h000;
            5158: color = 12'h000;
            5159: color = 12'h000;
            5160: color = 12'h000;
            5161: color = 12'h000;
            5162: color = 12'h000;
            5163: color = 12'h000;
            5164: color = 12'h000;
            5165: color = 12'h000;
            5166: color = 12'h000;
            5167: color = 12'h000;
            5168: color = 12'h000;
            5169: color = 12'h888;
            5170: color = 12'hFFF;
            5171: color = 12'hFFF;
            5172: color = 12'hFFF;
            5173: color = 12'hFFF;
            5174: color = 12'hFFF;
            5175: color = 12'hFFF;
            5176: color = 12'hFFF;
            5177: color = 12'hFFF;
            5178: color = 12'hFFF;
            5179: color = 12'hFFF;
            5180: color = 12'hFFF;
            5181: color = 12'h777;
            5182: color = 12'h000;
            5183: color = 12'h000;
            5184: color = 12'h000;
            5185: color = 12'h000;
            5186: color = 12'h000;
            5187: color = 12'h000;
            5188: color = 12'h000;
            5189: color = 12'h000;
            5190: color = 12'h000;
            5191: color = 12'h000;
            5192: color = 12'h000;
            5193: color = 12'h000;
            5194: color = 12'h000;
            5195: color = 12'h000;
            5196: color = 12'h000;
            5197: color = 12'h000;
            5198: color = 12'h000;
            5199: color = 12'h000;
            5200: color = 12'h000;
            5201: color = 12'h000;
            5202: color = 12'h000;
            5203: color = 12'h000;
            5204: color = 12'h000;
            5205: color = 12'h000;
            5206: color = 12'h000;
            5207: color = 12'h000;
            5208: color = 12'h000;
            5209: color = 12'h000;
            5210: color = 12'h000;
            5211: color = 12'h000;
            5212: color = 12'h000;
            5213: color = 12'h000;
            5214: color = 12'h000;
            5215: color = 12'h000;
            5216: color = 12'h000;
            5217: color = 12'h000;
            5218: color = 12'h000;
            5219: color = 12'h000;
            5220: color = 12'h000;
            5221: color = 12'h000;
            5222: color = 12'h000;
            5223: color = 12'h000;
            5224: color = 12'h000;
            5225: color = 12'h000;
            5226: color = 12'h000;
            5227: color = 12'h000;
            5228: color = 12'h000;
            5229: color = 12'h000;
            5230: color = 12'h000;
            5231: color = 12'h000;
            5232: color = 12'h000;
            5233: color = 12'h000;
            5234: color = 12'h000;
            5235: color = 12'h000;
            5236: color = 12'h000;
            5237: color = 12'h000;
            5238: color = 12'h000;
            5239: color = 12'h000;
            5240: color = 12'h000;
            5241: color = 12'h000;
            5242: color = 12'h000;
            5243: color = 12'hFFF;
            5244: color = 12'hFFF;
            5245: color = 12'hFFF;
            5246: color = 12'hFFF;
            5247: color = 12'hFFF;
            5248: color = 12'hFFF;
            5249: color = 12'hFFF;
            5250: color = 12'hFFF;
            5251: color = 12'hFFF;
            5252: color = 12'hFFF;
            5253: color = 12'hFFF;
            5254: color = 12'hFFF;
            5255: color = 12'hFFF;
            5256: color = 12'hFFF;
            5257: color = 12'hFFF;
            5258: color = 12'h000;
            5259: color = 12'h000;
            5260: color = 12'h000;
            5261: color = 12'h000;
            5262: color = 12'h000;
            5263: color = 12'h000;
            5264: color = 12'h000;
            5265: color = 12'h000;
            5266: color = 12'h000;
            5267: color = 12'h000;
            5268: color = 12'h000;
            5269: color = 12'h000;
            5270: color = 12'h000;
            5271: color = 12'h000;
            5272: color = 12'h000;
            5273: color = 12'h000;
            5274: color = 12'h000;
            5275: color = 12'h000;
            5276: color = 12'h777;
            5277: color = 12'h888;
            5278: color = 12'h777;
            5279: color = 12'h000;
            5280: color = 12'h000;
            5281: color = 12'h000;
            5282: color = 12'h000;
            5283: color = 12'h000;
            5284: color = 12'h000;
            5285: color = 12'h000;
            5286: color = 12'h000;
            5287: color = 12'h000;
            5288: color = 12'h000;
            5289: color = 12'h000;
            5290: color = 12'h000;
            5291: color = 12'h000;
            5292: color = 12'h000;
            5293: color = 12'h000;
            5294: color = 12'h000;
            5295: color = 12'h000;
            5296: color = 12'h000;
            5297: color = 12'h000;
            5298: color = 12'h000;
            5299: color = 12'h000;
            5300: color = 12'h000;
            5301: color = 12'h000;
            5302: color = 12'h000;
            5303: color = 12'h000;
            5304: color = 12'h000;
            5305: color = 12'h000;
            5306: color = 12'h000;
            5307: color = 12'h000;
            5308: color = 12'h000;
            5309: color = 12'h000;
            5310: color = 12'h000;
            5311: color = 12'h000;
            5312: color = 12'h000;
            5313: color = 12'h000;
            5314: color = 12'h000;
            5315: color = 12'h000;
            5316: color = 12'h000;
            5317: color = 12'h000;
            5318: color = 12'h777;
            5319: color = 12'h888;
            5320: color = 12'h777;
            5321: color = 12'h000;
            5322: color = 12'h000;
            5323: color = 12'h000;
            5324: color = 12'h000;
            5325: color = 12'h000;
            5326: color = 12'h000;
            5327: color = 12'h000;
            5328: color = 12'h000;
            5329: color = 12'h000;
            5330: color = 12'h000;
            5331: color = 12'h000;
            5332: color = 12'h000;
            5333: color = 12'h000;
            5334: color = 12'h000;
            5335: color = 12'h000;
            5336: color = 12'h000;
            5337: color = 12'h000;
            5338: color = 12'h000;
            5339: color = 12'h000;
            5340: color = 12'h000;
            5341: color = 12'h000;
            5342: color = 12'h000;
            5343: color = 12'h000;
            5344: color = 12'h000;
            5345: color = 12'h000;
            5346: color = 12'h000;
            5347: color = 12'h000;
            5348: color = 12'h000;
            5349: color = 12'h888;
            5350: color = 12'hFFF;
            5351: color = 12'hFFF;
            5352: color = 12'hFFF;
            5353: color = 12'hFFF;
            5354: color = 12'hFFF;
            5355: color = 12'hFFF;
            5356: color = 12'hFFF;
            5357: color = 12'hFFF;
            5358: color = 12'hFFF;
            5359: color = 12'hFFF;
            5360: color = 12'h000;
            5361: color = 12'h000;
            5362: color = 12'h000;
            5363: color = 12'h777;
            5364: color = 12'h888;
            5365: color = 12'h777;
            5366: color = 12'h000;
            5367: color = 12'h000;
            5368: color = 12'h000;
            5369: color = 12'h000;
            5370: color = 12'h000;
            5371: color = 12'h000;
            5372: color = 12'h000;
            5373: color = 12'h000;
            5374: color = 12'h000;
            5375: color = 12'h000;
            5376: color = 12'h000;
            5377: color = 12'h000;
            5378: color = 12'h000;
            5379: color = 12'h000;
            5380: color = 12'h000;
            5381: color = 12'h000;
            5382: color = 12'h000;
            5383: color = 12'h000;
            5384: color = 12'h000;
            5385: color = 12'h000;
            5386: color = 12'h000;
            5387: color = 12'h000;
            5388: color = 12'h000;
            5389: color = 12'h000;
            5390: color = 12'h000;
            5391: color = 12'h000;
            5392: color = 12'h000;
            5393: color = 12'h000;
            5394: color = 12'h000;
            5395: color = 12'h000;
            5396: color = 12'h000;
            5397: color = 12'h000;
            5398: color = 12'h000;
            5399: color = 12'h777;
            5400: color = 12'h888;
            5401: color = 12'h777;
            5402: color = 12'h000;
            5403: color = 12'h000;
            5404: color = 12'h000;
            5405: color = 12'h000;
            5406: color = 12'h000;
            5407: color = 12'h000;
            5408: color = 12'h000;
            5409: color = 12'h000;
            5410: color = 12'h000;
            5411: color = 12'h000;
            5412: color = 12'h000;
            5413: color = 12'h000;
            5414: color = 12'h000;
            5415: color = 12'h000;
            5416: color = 12'h000;
            5417: color = 12'h000;
            5418: color = 12'h000;
            5419: color = 12'h000;
            5420: color = 12'h000;
            5421: color = 12'h000;
            5422: color = 12'h000;
            5423: color = 12'h000;
            5424: color = 12'h000;
            5425: color = 12'h000;
            5426: color = 12'h000;
            5427: color = 12'h000;
            5428: color = 12'h000;
            5429: color = 12'h000;
            5430: color = 12'h000;
            5431: color = 12'h000;
            5432: color = 12'h000;
            5433: color = 12'h000;
            5434: color = 12'h000;
            5435: color = 12'h000;
            5436: color = 12'h000;
            5437: color = 12'h000;
            5438: color = 12'h000;
            5439: color = 12'h000;
            5440: color = 12'h000;
            5441: color = 12'h000;
            5442: color = 12'h000;
            5443: color = 12'h000;
            5444: color = 12'h000;
            5445: color = 12'h000;
            5446: color = 12'h000;
            5447: color = 12'h000;
            5448: color = 12'h000;
            5449: color = 12'h000;
            5450: color = 12'h000;
            5451: color = 12'h000;
            5452: color = 12'h000;
            5453: color = 12'h000;
            5454: color = 12'h000;
            5455: color = 12'h000;
            5456: color = 12'h000;
            5457: color = 12'h000;
            5458: color = 12'h000;
            5459: color = 12'h000;
            5460: color = 12'h000;
            5461: color = 12'h000;
            5462: color = 12'h000;
            5463: color = 12'h000;
            5464: color = 12'h000;
            5465: color = 12'h000;
            5466: color = 12'h000;
            5467: color = 12'h000;
            5468: color = 12'h000;
            5469: color = 12'h000;
            5470: color = 12'h000;
            5471: color = 12'h000;
            5472: color = 12'h000;
            5473: color = 12'h000;
            5474: color = 12'h000;
            5475: color = 12'h000;
            5476: color = 12'h000;
            5477: color = 12'h000;
            5478: color = 12'h000;
            5479: color = 12'h000;
            5480: color = 12'h000;
            5481: color = 12'h000;
            5482: color = 12'h000;
            5483: color = 12'h000;
            5484: color = 12'h000;
            5485: color = 12'h000;
            5486: color = 12'h000;
            5487: color = 12'h000;
            5488: color = 12'h000;
            5489: color = 12'h888;
            5490: color = 12'hFFF;
            5491: color = 12'hFFF;
            5492: color = 12'hFFF;
            5493: color = 12'hFFF;
            5494: color = 12'hFFF;
            5495: color = 12'hFFF;
            5496: color = 12'hFFF;
            5497: color = 12'hFFF;
            5498: color = 12'hFFF;
            5499: color = 12'hFFF;
            5500: color = 12'hFFF;
            5501: color = 12'h888;
            5502: color = 12'h000;
            5503: color = 12'h000;
            5504: color = 12'h000;
            5505: color = 12'h000;
            5506: color = 12'h000;
            5507: color = 12'h000;
            5508: color = 12'h000;
            5509: color = 12'h000;
            5510: color = 12'h000;
            5511: color = 12'h000;
            5512: color = 12'h000;
            5513: color = 12'h000;
            5514: color = 12'h000;
            5515: color = 12'h000;
            5516: color = 12'h000;
            5517: color = 12'h000;
            5518: color = 12'h000;
            5519: color = 12'h000;
            5520: color = 12'h000;
            5521: color = 12'h000;
            5522: color = 12'h000;
            5523: color = 12'h000;
            5524: color = 12'h000;
            5525: color = 12'h000;
            5526: color = 12'h000;
            5527: color = 12'h000;
            5528: color = 12'h000;
            5529: color = 12'h000;
            5530: color = 12'h000;
            5531: color = 12'h000;
            5532: color = 12'h000;
            5533: color = 12'h000;
            5534: color = 12'h000;
            5535: color = 12'h000;
            5536: color = 12'h000;
            5537: color = 12'h000;
            5538: color = 12'h000;
            5539: color = 12'h000;
            5540: color = 12'h000;
            5541: color = 12'h000;
            5542: color = 12'h000;
            5543: color = 12'h000;
            5544: color = 12'h000;
            5545: color = 12'h000;
            5546: color = 12'h000;
            5547: color = 12'h000;
            5548: color = 12'h000;
            5549: color = 12'h000;
            5550: color = 12'h000;
            5551: color = 12'h000;
            5552: color = 12'h000;
            5553: color = 12'h000;
            5554: color = 12'h000;
            5555: color = 12'h000;
            5556: color = 12'h000;
            5557: color = 12'h000;
            5558: color = 12'h000;
            5559: color = 12'h000;
            5560: color = 12'h000;
            5561: color = 12'h000;
            5562: color = 12'h000;
            5563: color = 12'hFFF;
            5564: color = 12'hFFF;
            5565: color = 12'hFFF;
            5566: color = 12'hFFF;
            5567: color = 12'hFFF;
            5568: color = 12'hFFF;
            5569: color = 12'hFFF;
            5570: color = 12'hFFF;
            5571: color = 12'hFFF;
            5572: color = 12'hFFF;
            5573: color = 12'hFFF;
            5574: color = 12'hFFF;
            5575: color = 12'hFFF;
            5576: color = 12'hFFF;
            5577: color = 12'hEEE;
            5578: color = 12'h000;
            5579: color = 12'h000;
            5580: color = 12'h000;
            5581: color = 12'h000;
            5582: color = 12'h000;
            5583: color = 12'h000;
            5584: color = 12'h000;
            5585: color = 12'h000;
            5586: color = 12'h000;
            5587: color = 12'h000;
            5588: color = 12'h000;
            5589: color = 12'h000;
            5590: color = 12'h000;
            5591: color = 12'h000;
            5592: color = 12'h000;
            5593: color = 12'h000;
            5594: color = 12'h000;
            5595: color = 12'h000;
            5596: color = 12'hFFF;
            5597: color = 12'hFFF;
            5598: color = 12'hFFF;
            5599: color = 12'h000;
            5600: color = 12'h000;
            5601: color = 12'h000;
            5602: color = 12'h000;
            5603: color = 12'h000;
            5604: color = 12'h000;
            5605: color = 12'h000;
            5606: color = 12'h000;
            5607: color = 12'h000;
            5608: color = 12'h000;
            5609: color = 12'h000;
            5610: color = 12'h000;
            5611: color = 12'h000;
            5612: color = 12'h000;
            5613: color = 12'h000;
            5614: color = 12'h000;
            5615: color = 12'h000;
            5616: color = 12'h000;
            5617: color = 12'h000;
            5618: color = 12'h000;
            5619: color = 12'h000;
            5620: color = 12'h000;
            5621: color = 12'h000;
            5622: color = 12'h000;
            5623: color = 12'h000;
            5624: color = 12'h000;
            5625: color = 12'h000;
            5626: color = 12'h000;
            5627: color = 12'h000;
            5628: color = 12'h000;
            5629: color = 12'h000;
            5630: color = 12'h000;
            5631: color = 12'h000;
            5632: color = 12'h000;
            5633: color = 12'h000;
            5634: color = 12'h000;
            5635: color = 12'h000;
            5636: color = 12'h000;
            5637: color = 12'h000;
            5638: color = 12'hFFF;
            5639: color = 12'hFFF;
            5640: color = 12'hFFF;
            5641: color = 12'h000;
            5642: color = 12'h000;
            5643: color = 12'h000;
            5644: color = 12'h000;
            5645: color = 12'h000;
            5646: color = 12'h000;
            5647: color = 12'h000;
            5648: color = 12'h000;
            5649: color = 12'h000;
            5650: color = 12'h000;
            5651: color = 12'h000;
            5652: color = 12'h000;
            5653: color = 12'h000;
            5654: color = 12'h000;
            5655: color = 12'h000;
            5656: color = 12'h000;
            5657: color = 12'h000;
            5658: color = 12'h000;
            5659: color = 12'h000;
            5660: color = 12'h000;
            5661: color = 12'h000;
            5662: color = 12'h000;
            5663: color = 12'h000;
            5664: color = 12'h000;
            5665: color = 12'h000;
            5666: color = 12'h000;
            5667: color = 12'h000;
            5668: color = 12'h000;
            5669: color = 12'h888;
            5670: color = 12'hFFF;
            5671: color = 12'hFFF;
            5672: color = 12'hFFF;
            5673: color = 12'hFFF;
            5674: color = 12'hFFF;
            5675: color = 12'hFFF;
            5676: color = 12'hFFF;
            5677: color = 12'hFFF;
            5678: color = 12'hFFF;
            5679: color = 12'hEEE;
            5680: color = 12'h000;
            5681: color = 12'h000;
            5682: color = 12'h000;
            5683: color = 12'hFFF;
            5684: color = 12'hFFF;
            5685: color = 12'hFFF;
            5686: color = 12'h000;
            5687: color = 12'h000;
            5688: color = 12'h000;
            5689: color = 12'h000;
            5690: color = 12'h000;
            5691: color = 12'h000;
            5692: color = 12'h000;
            5693: color = 12'h000;
            5694: color = 12'h000;
            5695: color = 12'h000;
            5696: color = 12'h000;
            5697: color = 12'h000;
            5698: color = 12'h000;
            5699: color = 12'h000;
            5700: color = 12'h000;
            5701: color = 12'h000;
            5702: color = 12'h000;
            5703: color = 12'h000;
            5704: color = 12'h000;
            5705: color = 12'h000;
            5706: color = 12'h000;
            5707: color = 12'h000;
            5708: color = 12'h000;
            5709: color = 12'h000;
            5710: color = 12'h000;
            5711: color = 12'h000;
            5712: color = 12'h000;
            5713: color = 12'h000;
            5714: color = 12'h000;
            5715: color = 12'h000;
            5716: color = 12'h000;
            5717: color = 12'h000;
            5718: color = 12'h000;
            5719: color = 12'hFFF;
            5720: color = 12'hFFF;
            5721: color = 12'hFFF;
            5722: color = 12'h000;
            5723: color = 12'h000;
            5724: color = 12'h000;
            5725: color = 12'h000;
            5726: color = 12'h000;
            5727: color = 12'h000;
            5728: color = 12'h000;
            5729: color = 12'h000;
            5730: color = 12'h000;
            5731: color = 12'h000;
            5732: color = 12'h000;
            5733: color = 12'h000;
            5734: color = 12'h000;
            5735: color = 12'h000;
            5736: color = 12'h000;
            5737: color = 12'h000;
            5738: color = 12'h000;
            5739: color = 12'h000;
            5740: color = 12'h000;
            5741: color = 12'h000;
            5742: color = 12'h000;
            5743: color = 12'h000;
            5744: color = 12'h000;
            5745: color = 12'h000;
            5746: color = 12'h000;
            5747: color = 12'h000;
            5748: color = 12'h000;
            5749: color = 12'h000;
            5750: color = 12'h000;
            5751: color = 12'h000;
            5752: color = 12'h000;
            5753: color = 12'h000;
            5754: color = 12'h000;
            5755: color = 12'h000;
            5756: color = 12'h000;
            5757: color = 12'h000;
            5758: color = 12'h000;
            5759: color = 12'h000;
            5760: color = 12'h000;
            5761: color = 12'h000;
            5762: color = 12'h000;
            5763: color = 12'h000;
            5764: color = 12'h000;
            5765: color = 12'h000;
            5766: color = 12'h000;
            5767: color = 12'h000;
            5768: color = 12'h000;
            5769: color = 12'h000;
            5770: color = 12'h000;
            5771: color = 12'h000;
            5772: color = 12'h000;
            5773: color = 12'h000;
            5774: color = 12'h000;
            5775: color = 12'h000;
            5776: color = 12'h000;
            5777: color = 12'h000;
            5778: color = 12'h000;
            5779: color = 12'h000;
            5780: color = 12'h000;
            5781: color = 12'h000;
            5782: color = 12'h000;
            5783: color = 12'h000;
            5784: color = 12'h000;
            5785: color = 12'h000;
            5786: color = 12'h000;
            5787: color = 12'h000;
            5788: color = 12'h000;
            5789: color = 12'h000;
            5790: color = 12'h000;
            5791: color = 12'h000;
            5792: color = 12'h000;
            5793: color = 12'h000;
            5794: color = 12'h000;
            5795: color = 12'h000;
            5796: color = 12'h000;
            5797: color = 12'h000;
            5798: color = 12'h000;
            5799: color = 12'h000;
            5800: color = 12'h000;
            5801: color = 12'h000;
            5802: color = 12'h000;
            5803: color = 12'h000;
            5804: color = 12'h000;
            5805: color = 12'h000;
            5806: color = 12'h000;
            5807: color = 12'h000;
            5808: color = 12'h000;
            5809: color = 12'h888;
            5810: color = 12'hFFF;
            5811: color = 12'hFFF;
            5812: color = 12'h888;
            5813: color = 12'h000;
            5814: color = 12'h000;
            5815: color = 12'h000;
            5816: color = 12'h000;
            5817: color = 12'h000;
            5818: color = 12'h000;
            5819: color = 12'h000;
            5820: color = 12'h000;
            5821: color = 12'h888;
            5822: color = 12'hFFF;
            5823: color = 12'hFFF;
            5824: color = 12'h777;
            5825: color = 12'h000;
            5826: color = 12'h000;
            5827: color = 12'h000;
            5828: color = 12'h000;
            5829: color = 12'h000;
            5830: color = 12'h000;
            5831: color = 12'h000;
            5832: color = 12'h000;
            5833: color = 12'h000;
            5834: color = 12'h000;
            5835: color = 12'h000;
            5836: color = 12'h000;
            5837: color = 12'h000;
            5838: color = 12'h000;
            5839: color = 12'h000;
            5840: color = 12'h000;
            5841: color = 12'h000;
            5842: color = 12'h000;
            5843: color = 12'h000;
            5844: color = 12'h000;
            5845: color = 12'h000;
            5846: color = 12'h000;
            5847: color = 12'h000;
            5848: color = 12'h000;
            5849: color = 12'h000;
            5850: color = 12'h000;
            5851: color = 12'h000;
            5852: color = 12'h000;
            5853: color = 12'h000;
            5854: color = 12'h777;
            5855: color = 12'hFFF;
            5856: color = 12'hFFF;
            5857: color = 12'hFFF;
            5858: color = 12'hFFF;
            5859: color = 12'hFFF;
            5860: color = 12'hFFF;
            5861: color = 12'hEEE;
            5862: color = 12'h000;
            5863: color = 12'h000;
            5864: color = 12'h000;
            5865: color = 12'h000;
            5866: color = 12'h777;
            5867: color = 12'hFFF;
            5868: color = 12'hFFF;
            5869: color = 12'hFFF;
            5870: color = 12'hFFF;
            5871: color = 12'hFFF;
            5872: color = 12'hFFF;
            5873: color = 12'hEEE;
            5874: color = 12'h000;
            5875: color = 12'h000;
            5876: color = 12'h000;
            5877: color = 12'h000;
            5878: color = 12'h000;
            5879: color = 12'h000;
            5880: color = 12'h000;
            5881: color = 12'h000;
            5882: color = 12'h000;
            5883: color = 12'hFFF;
            5884: color = 12'hFFF;
            5885: color = 12'hFFF;
            5886: color = 12'h111;
            5887: color = 12'h000;
            5888: color = 12'h000;
            5889: color = 12'h000;
            5890: color = 12'h000;
            5891: color = 12'h000;
            5892: color = 12'h000;
            5893: color = 12'h000;
            5894: color = 12'h000;
            5895: color = 12'h000;
            5896: color = 12'h000;
            5897: color = 12'h000;
            5898: color = 12'h000;
            5899: color = 12'h000;
            5900: color = 12'h000;
            5901: color = 12'h000;
            5902: color = 12'h000;
            5903: color = 12'h000;
            5904: color = 12'h000;
            5905: color = 12'h000;
            5906: color = 12'h000;
            5907: color = 12'h000;
            5908: color = 12'h000;
            5909: color = 12'h000;
            5910: color = 12'h000;
            5911: color = 12'h000;
            5912: color = 12'h000;
            5913: color = 12'h000;
            5914: color = 12'h000;
            5915: color = 12'h000;
            5916: color = 12'hFFF;
            5917: color = 12'hFFF;
            5918: color = 12'hFFF;
            5919: color = 12'h000;
            5920: color = 12'h000;
            5921: color = 12'h000;
            5922: color = 12'h000;
            5923: color = 12'h000;
            5924: color = 12'h000;
            5925: color = 12'h000;
            5926: color = 12'h000;
            5927: color = 12'h000;
            5928: color = 12'h000;
            5929: color = 12'h000;
            5930: color = 12'h000;
            5931: color = 12'h000;
            5932: color = 12'h000;
            5933: color = 12'h000;
            5934: color = 12'h000;
            5935: color = 12'h000;
            5936: color = 12'h000;
            5937: color = 12'h000;
            5938: color = 12'h000;
            5939: color = 12'h000;
            5940: color = 12'h000;
            5941: color = 12'h000;
            5942: color = 12'h000;
            5943: color = 12'h000;
            5944: color = 12'h000;
            5945: color = 12'h000;
            5946: color = 12'h000;
            5947: color = 12'h000;
            5948: color = 12'h000;
            5949: color = 12'h000;
            5950: color = 12'h000;
            5951: color = 12'h000;
            5952: color = 12'h000;
            5953: color = 12'h000;
            5954: color = 12'h000;
            5955: color = 12'h000;
            5956: color = 12'h000;
            5957: color = 12'h000;
            5958: color = 12'hFFF;
            5959: color = 12'hFFF;
            5960: color = 12'hFFF;
            5961: color = 12'h000;
            5962: color = 12'h000;
            5963: color = 12'h000;
            5964: color = 12'h000;
            5965: color = 12'h000;
            5966: color = 12'h000;
            5967: color = 12'h000;
            5968: color = 12'h000;
            5969: color = 12'h000;
            5970: color = 12'h000;
            5971: color = 12'h000;
            5972: color = 12'h000;
            5973: color = 12'h000;
            5974: color = 12'h000;
            5975: color = 12'h000;
            5976: color = 12'h000;
            5977: color = 12'h000;
            5978: color = 12'h000;
            5979: color = 12'h000;
            5980: color = 12'h000;
            5981: color = 12'h000;
            5982: color = 12'h000;
            5983: color = 12'h000;
            5984: color = 12'h000;
            5985: color = 12'h000;
            5986: color = 12'h777;
            5987: color = 12'hFFF;
            5988: color = 12'hFFF;
            5989: color = 12'h888;
            5990: color = 12'h000;
            5991: color = 12'h000;
            5992: color = 12'h000;
            5993: color = 12'h000;
            5994: color = 12'h000;
            5995: color = 12'h000;
            5996: color = 12'h000;
            5997: color = 12'h000;
            5998: color = 12'h000;
            5999: color = 12'h000;
            6000: color = 12'h000;
            6001: color = 12'h000;
            6002: color = 12'h000;
            6003: color = 12'hFFF;
            6004: color = 12'hFFF;
            6005: color = 12'hFFF;
            6006: color = 12'h000;
            6007: color = 12'h000;
            6008: color = 12'h000;
            6009: color = 12'h000;
            6010: color = 12'h000;
            6011: color = 12'h000;
            6012: color = 12'h000;
            6013: color = 12'h000;
            6014: color = 12'h000;
            6015: color = 12'h000;
            6016: color = 12'h000;
            6017: color = 12'h000;
            6018: color = 12'h000;
            6019: color = 12'h000;
            6020: color = 12'h000;
            6021: color = 12'h000;
            6022: color = 12'h000;
            6023: color = 12'h000;
            6024: color = 12'h000;
            6025: color = 12'h000;
            6026: color = 12'h000;
            6027: color = 12'h000;
            6028: color = 12'h000;
            6029: color = 12'h000;
            6030: color = 12'h000;
            6031: color = 12'h000;
            6032: color = 12'h000;
            6033: color = 12'h000;
            6034: color = 12'h000;
            6035: color = 12'h000;
            6036: color = 12'h000;
            6037: color = 12'h000;
            6038: color = 12'h000;
            6039: color = 12'hFFF;
            6040: color = 12'hFFF;
            6041: color = 12'hFFF;
            6042: color = 12'h000;
            6043: color = 12'h000;
            6044: color = 12'h000;
            6045: color = 12'h000;
            6046: color = 12'h000;
            6047: color = 12'h000;
            6048: color = 12'h000;
            6049: color = 12'h000;
            6050: color = 12'h000;
            6051: color = 12'h000;
            6052: color = 12'h000;
            6053: color = 12'h000;
            6054: color = 12'h000;
            6055: color = 12'h000;
            6056: color = 12'h000;
            6057: color = 12'h000;
            6058: color = 12'h000;
            6059: color = 12'h000;
            6060: color = 12'h000;
            6061: color = 12'h000;
            6062: color = 12'h000;
            6063: color = 12'h000;
            6064: color = 12'h000;
            6065: color = 12'h000;
            6066: color = 12'h000;
            6067: color = 12'h000;
            6068: color = 12'h000;
            6069: color = 12'h000;
            6070: color = 12'h000;
            6071: color = 12'h000;
            6072: color = 12'h000;
            6073: color = 12'h000;
            6074: color = 12'h000;
            6075: color = 12'h000;
            6076: color = 12'h000;
            6077: color = 12'h000;
            6078: color = 12'h000;
            6079: color = 12'h000;
            6080: color = 12'h000;
            6081: color = 12'h000;
            6082: color = 12'h000;
            6083: color = 12'h000;
            6084: color = 12'h000;
            6085: color = 12'h000;
            6086: color = 12'h000;
            6087: color = 12'h000;
            6088: color = 12'h000;
            6089: color = 12'h000;
            6090: color = 12'h000;
            6091: color = 12'h000;
            6092: color = 12'h000;
            6093: color = 12'h000;
            6094: color = 12'h000;
            6095: color = 12'h000;
            6096: color = 12'h000;
            6097: color = 12'h000;
            6098: color = 12'h000;
            6099: color = 12'h000;
            6100: color = 12'h000;
            6101: color = 12'h000;
            6102: color = 12'h000;
            6103: color = 12'h000;
            6104: color = 12'h000;
            6105: color = 12'h000;
            6106: color = 12'h000;
            6107: color = 12'h000;
            6108: color = 12'h000;
            6109: color = 12'h000;
            6110: color = 12'h000;
            6111: color = 12'h000;
            6112: color = 12'h000;
            6113: color = 12'h000;
            6114: color = 12'h000;
            6115: color = 12'h000;
            6116: color = 12'h000;
            6117: color = 12'h000;
            6118: color = 12'h000;
            6119: color = 12'h000;
            6120: color = 12'h000;
            6121: color = 12'h000;
            6122: color = 12'h000;
            6123: color = 12'h000;
            6124: color = 12'h000;
            6125: color = 12'h000;
            6126: color = 12'h000;
            6127: color = 12'h000;
            6128: color = 12'h000;
            6129: color = 12'h888;
            6130: color = 12'hFFF;
            6131: color = 12'hFFF;
            6132: color = 12'h777;
            6133: color = 12'h000;
            6134: color = 12'h000;
            6135: color = 12'h000;
            6136: color = 12'h000;
            6137: color = 12'h000;
            6138: color = 12'h000;
            6139: color = 12'h000;
            6140: color = 12'h000;
            6141: color = 12'h888;
            6142: color = 12'hFFF;
            6143: color = 12'hFFF;
            6144: color = 12'h777;
            6145: color = 12'h000;
            6146: color = 12'h777;
            6147: color = 12'h888;
            6148: color = 12'h777;
            6149: color = 12'h000;
            6150: color = 12'h444;
            6151: color = 12'h888;
            6152: color = 12'h888;
            6153: color = 12'h888;
            6154: color = 12'h777;
            6155: color = 12'h000;
            6156: color = 12'h000;
            6157: color = 12'h000;
            6158: color = 12'h000;
            6159: color = 12'h000;
            6160: color = 12'h000;
            6161: color = 12'h777;
            6162: color = 12'h888;
            6163: color = 12'h888;
            6164: color = 12'h888;
            6165: color = 12'h888;
            6166: color = 12'h888;
            6167: color = 12'h888;
            6168: color = 12'h888;
            6169: color = 12'h777;
            6170: color = 12'h000;
            6171: color = 12'h000;
            6172: color = 12'h000;
            6173: color = 12'h000;
            6174: color = 12'h888;
            6175: color = 12'hFFF;
            6176: color = 12'hFFF;
            6177: color = 12'hFFF;
            6178: color = 12'hFFF;
            6179: color = 12'hFFF;
            6180: color = 12'hFFF;
            6181: color = 12'hFFF;
            6182: color = 12'h000;
            6183: color = 12'h000;
            6184: color = 12'h000;
            6185: color = 12'h000;
            6186: color = 12'h888;
            6187: color = 12'hFFF;
            6188: color = 12'hFFF;
            6189: color = 12'hFFF;
            6190: color = 12'hFFF;
            6191: color = 12'hFFF;
            6192: color = 12'hFFF;
            6193: color = 12'hFFF;
            6194: color = 12'h000;
            6195: color = 12'h000;
            6196: color = 12'h000;
            6197: color = 12'h000;
            6198: color = 12'h000;
            6199: color = 12'h000;
            6200: color = 12'h000;
            6201: color = 12'h000;
            6202: color = 12'h000;
            6203: color = 12'hFFF;
            6204: color = 12'hFFF;
            6205: color = 12'hFFF;
            6206: color = 12'h000;
            6207: color = 12'h000;
            6208: color = 12'h000;
            6209: color = 12'h000;
            6210: color = 12'h000;
            6211: color = 12'h000;
            6212: color = 12'h000;
            6213: color = 12'h000;
            6214: color = 12'h000;
            6215: color = 12'h000;
            6216: color = 12'h000;
            6217: color = 12'h000;
            6218: color = 12'h000;
            6219: color = 12'h444;
            6220: color = 12'h888;
            6221: color = 12'h888;
            6222: color = 12'h888;
            6223: color = 12'h888;
            6224: color = 12'h888;
            6225: color = 12'h888;
            6226: color = 12'h888;
            6227: color = 12'h888;
            6228: color = 12'h888;
            6229: color = 12'h777;
            6230: color = 12'h000;
            6231: color = 12'h000;
            6232: color = 12'h000;
            6233: color = 12'h000;
            6234: color = 12'h444;
            6235: color = 12'h888;
            6236: color = 12'hFFF;
            6237: color = 12'hFFF;
            6238: color = 12'hFFF;
            6239: color = 12'h888;
            6240: color = 12'h444;
            6241: color = 12'h000;
            6242: color = 12'h000;
            6243: color = 12'h000;
            6244: color = 12'h000;
            6245: color = 12'h000;
            6246: color = 12'h444;
            6247: color = 12'h888;
            6248: color = 12'h888;
            6249: color = 12'h888;
            6250: color = 12'h888;
            6251: color = 12'h888;
            6252: color = 12'h888;
            6253: color = 12'h888;
            6254: color = 12'h888;
            6255: color = 12'h444;
            6256: color = 12'h000;
            6257: color = 12'h777;
            6258: color = 12'h888;
            6259: color = 12'h777;
            6260: color = 12'h000;
            6261: color = 12'h444;
            6262: color = 12'h888;
            6263: color = 12'h888;
            6264: color = 12'h888;
            6265: color = 12'h777;
            6266: color = 12'h000;
            6267: color = 12'h000;
            6268: color = 12'h000;
            6269: color = 12'h000;
            6270: color = 12'h000;
            6271: color = 12'h000;
            6272: color = 12'h000;
            6273: color = 12'h000;
            6274: color = 12'h000;
            6275: color = 12'h000;
            6276: color = 12'h444;
            6277: color = 12'h888;
            6278: color = 12'hFFF;
            6279: color = 12'hFFF;
            6280: color = 12'hFFF;
            6281: color = 12'h888;
            6282: color = 12'h444;
            6283: color = 12'h000;
            6284: color = 12'h000;
            6285: color = 12'h000;
            6286: color = 12'h000;
            6287: color = 12'h000;
            6288: color = 12'h444;
            6289: color = 12'h888;
            6290: color = 12'h888;
            6291: color = 12'h888;
            6292: color = 12'h888;
            6293: color = 12'h888;
            6294: color = 12'h444;
            6295: color = 12'h000;
            6296: color = 12'h000;
            6297: color = 12'h000;
            6298: color = 12'h000;
            6299: color = 12'h000;
            6300: color = 12'h000;
            6301: color = 12'h000;
            6302: color = 12'h000;
            6303: color = 12'h000;
            6304: color = 12'h000;
            6305: color = 12'h000;
            6306: color = 12'h888;
            6307: color = 12'hFFF;
            6308: color = 12'hFFF;
            6309: color = 12'h777;
            6310: color = 12'h000;
            6311: color = 12'h000;
            6312: color = 12'h000;
            6313: color = 12'h000;
            6314: color = 12'h000;
            6315: color = 12'h000;
            6316: color = 12'h000;
            6317: color = 12'h000;
            6318: color = 12'h000;
            6319: color = 12'h000;
            6320: color = 12'h000;
            6321: color = 12'h444;
            6322: color = 12'h888;
            6323: color = 12'hFFF;
            6324: color = 12'hFFF;
            6325: color = 12'hFFF;
            6326: color = 12'h888;
            6327: color = 12'h444;
            6328: color = 12'h000;
            6329: color = 12'h000;
            6330: color = 12'h444;
            6331: color = 12'h888;
            6332: color = 12'h888;
            6333: color = 12'h888;
            6334: color = 12'h888;
            6335: color = 12'h888;
            6336: color = 12'h888;
            6337: color = 12'h888;
            6338: color = 12'h888;
            6339: color = 12'h888;
            6340: color = 12'h777;
            6341: color = 12'h000;
            6342: color = 12'h000;
            6343: color = 12'h000;
            6344: color = 12'h000;
            6345: color = 12'h444;
            6346: color = 12'h888;
            6347: color = 12'h888;
            6348: color = 12'h444;
            6349: color = 12'h000;
            6350: color = 12'h777;
            6351: color = 12'h888;
            6352: color = 12'h888;
            6353: color = 12'h888;
            6354: color = 12'h444;
            6355: color = 12'h000;
            6356: color = 12'h000;
            6357: color = 12'h444;
            6358: color = 12'h888;
            6359: color = 12'hFFF;
            6360: color = 12'hFFF;
            6361: color = 12'hFFF;
            6362: color = 12'h888;
            6363: color = 12'h444;
            6364: color = 12'h000;
            6365: color = 12'h000;
            6366: color = 12'h000;
            6367: color = 12'h000;
            6368: color = 12'h000;
            6369: color = 12'h000;
            6370: color = 12'h000;
            6371: color = 12'h000;
            6372: color = 12'h000;
            6373: color = 12'h000;
            6374: color = 12'h000;
            6375: color = 12'h000;
            6376: color = 12'h000;
            6377: color = 12'h000;
            6378: color = 12'h000;
            6379: color = 12'h000;
            6380: color = 12'h000;
            6381: color = 12'h000;
            6382: color = 12'h000;
            6383: color = 12'h000;
            6384: color = 12'h000;
            6385: color = 12'h000;
            6386: color = 12'h000;
            6387: color = 12'h000;
            6388: color = 12'h000;
            6389: color = 12'h000;
            6390: color = 12'h000;
            6391: color = 12'h000;
            6392: color = 12'h000;
            6393: color = 12'h000;
            6394: color = 12'h000;
            6395: color = 12'h000;
            6396: color = 12'h000;
            6397: color = 12'h000;
            6398: color = 12'h000;
            6399: color = 12'h000;
            6400: color = 12'h000;
            6401: color = 12'h000;
            6402: color = 12'h000;
            6403: color = 12'h000;
            6404: color = 12'h000;
            6405: color = 12'h000;
            6406: color = 12'h000;
            6407: color = 12'h000;
            6408: color = 12'h000;
            6409: color = 12'h000;
            6410: color = 12'h000;
            6411: color = 12'h000;
            6412: color = 12'h000;
            6413: color = 12'h000;
            6414: color = 12'h000;
            6415: color = 12'h000;
            6416: color = 12'h000;
            6417: color = 12'h000;
            6418: color = 12'h000;
            6419: color = 12'h000;
            6420: color = 12'h000;
            6421: color = 12'h000;
            6422: color = 12'h000;
            6423: color = 12'h000;
            6424: color = 12'h000;
            6425: color = 12'h000;
            6426: color = 12'h000;
            6427: color = 12'h000;
            6428: color = 12'h000;
            6429: color = 12'h000;
            6430: color = 12'h000;
            6431: color = 12'h000;
            6432: color = 12'h000;
            6433: color = 12'h000;
            6434: color = 12'h000;
            6435: color = 12'h000;
            6436: color = 12'h000;
            6437: color = 12'h000;
            6438: color = 12'h000;
            6439: color = 12'h000;
            6440: color = 12'h000;
            6441: color = 12'h000;
            6442: color = 12'h000;
            6443: color = 12'h000;
            6444: color = 12'h000;
            6445: color = 12'h000;
            6446: color = 12'h000;
            6447: color = 12'h000;
            6448: color = 12'h000;
            6449: color = 12'h888;
            6450: color = 12'hFFF;
            6451: color = 12'hFFF;
            6452: color = 12'h888;
            6453: color = 12'h000;
            6454: color = 12'h000;
            6455: color = 12'h000;
            6456: color = 12'h000;
            6457: color = 12'h000;
            6458: color = 12'h000;
            6459: color = 12'h000;
            6460: color = 12'h000;
            6461: color = 12'h888;
            6462: color = 12'hFFF;
            6463: color = 12'hFFF;
            6464: color = 12'h777;
            6465: color = 12'h000;
            6466: color = 12'hFFF;
            6467: color = 12'hFFF;
            6468: color = 12'hFFF;
            6469: color = 12'h111;
            6470: color = 12'h888;
            6471: color = 12'hFFF;
            6472: color = 12'hFFF;
            6473: color = 12'hFFF;
            6474: color = 12'hFFF;
            6475: color = 12'h111;
            6476: color = 12'h000;
            6477: color = 12'h000;
            6478: color = 12'h000;
            6479: color = 12'h000;
            6480: color = 12'h000;
            6481: color = 12'hFFF;
            6482: color = 12'hFFF;
            6483: color = 12'hFFF;
            6484: color = 12'hFFF;
            6485: color = 12'hFFF;
            6486: color = 12'hFFF;
            6487: color = 12'hFFF;
            6488: color = 12'hFFF;
            6489: color = 12'hFFF;
            6490: color = 12'h000;
            6491: color = 12'h000;
            6492: color = 12'h000;
            6493: color = 12'h000;
            6494: color = 12'h888;
            6495: color = 12'hFFF;
            6496: color = 12'hFFF;
            6497: color = 12'hFFF;
            6498: color = 12'hFFF;
            6499: color = 12'hFFF;
            6500: color = 12'hFFF;
            6501: color = 12'hEEE;
            6502: color = 12'h000;
            6503: color = 12'h000;
            6504: color = 12'h000;
            6505: color = 12'h000;
            6506: color = 12'h888;
            6507: color = 12'hFFF;
            6508: color = 12'hFFF;
            6509: color = 12'hFFF;
            6510: color = 12'hFFF;
            6511: color = 12'hFFF;
            6512: color = 12'hFFF;
            6513: color = 12'hEEE;
            6514: color = 12'h000;
            6515: color = 12'h000;
            6516: color = 12'h000;
            6517: color = 12'h000;
            6518: color = 12'h000;
            6519: color = 12'h000;
            6520: color = 12'h000;
            6521: color = 12'h000;
            6522: color = 12'h000;
            6523: color = 12'hFFF;
            6524: color = 12'hFFF;
            6525: color = 12'hFFF;
            6526: color = 12'h111;
            6527: color = 12'h000;
            6528: color = 12'h000;
            6529: color = 12'h000;
            6530: color = 12'h000;
            6531: color = 12'h000;
            6532: color = 12'h000;
            6533: color = 12'h000;
            6534: color = 12'h000;
            6535: color = 12'h000;
            6536: color = 12'h000;
            6537: color = 12'h000;
            6538: color = 12'h000;
            6539: color = 12'h888;
            6540: color = 12'hFFF;
            6541: color = 12'hFFF;
            6542: color = 12'hFFF;
            6543: color = 12'hFFF;
            6544: color = 12'hFFF;
            6545: color = 12'hFFF;
            6546: color = 12'hFFF;
            6547: color = 12'hFFF;
            6548: color = 12'hFFF;
            6549: color = 12'hFFF;
            6550: color = 12'h000;
            6551: color = 12'h000;
            6552: color = 12'h000;
            6553: color = 12'h000;
            6554: color = 12'h888;
            6555: color = 12'hFFF;
            6556: color = 12'hFFF;
            6557: color = 12'hFFF;
            6558: color = 12'hFFF;
            6559: color = 12'hFFF;
            6560: color = 12'h777;
            6561: color = 12'h000;
            6562: color = 12'h000;
            6563: color = 12'h000;
            6564: color = 12'h000;
            6565: color = 12'h000;
            6566: color = 12'h888;
            6567: color = 12'hFFF;
            6568: color = 12'hFFF;
            6569: color = 12'hFFF;
            6570: color = 12'hFFF;
            6571: color = 12'hFFF;
            6572: color = 12'hFFF;
            6573: color = 12'hFFF;
            6574: color = 12'hFFF;
            6575: color = 12'h777;
            6576: color = 12'h000;
            6577: color = 12'hFFF;
            6578: color = 12'hFFF;
            6579: color = 12'hFFF;
            6580: color = 12'h111;
            6581: color = 12'h888;
            6582: color = 12'hFFF;
            6583: color = 12'hFFF;
            6584: color = 12'hFFF;
            6585: color = 12'hFFF;
            6586: color = 12'h111;
            6587: color = 12'h000;
            6588: color = 12'h000;
            6589: color = 12'h000;
            6590: color = 12'h000;
            6591: color = 12'h000;
            6592: color = 12'h000;
            6593: color = 12'h000;
            6594: color = 12'h000;
            6595: color = 12'h000;
            6596: color = 12'h888;
            6597: color = 12'hFFF;
            6598: color = 12'hFFF;
            6599: color = 12'hFFF;
            6600: color = 12'hFFF;
            6601: color = 12'hFFF;
            6602: color = 12'h777;
            6603: color = 12'h000;
            6604: color = 12'h000;
            6605: color = 12'h000;
            6606: color = 12'h000;
            6607: color = 12'h000;
            6608: color = 12'h888;
            6609: color = 12'hFFF;
            6610: color = 12'hFFF;
            6611: color = 12'hFFF;
            6612: color = 12'hFFF;
            6613: color = 12'hFFF;
            6614: color = 12'h777;
            6615: color = 12'h000;
            6616: color = 12'h000;
            6617: color = 12'h000;
            6618: color = 12'h000;
            6619: color = 12'h000;
            6620: color = 12'h000;
            6621: color = 12'h000;
            6622: color = 12'h000;
            6623: color = 12'h000;
            6624: color = 12'h000;
            6625: color = 12'h000;
            6626: color = 12'h777;
            6627: color = 12'hFFF;
            6628: color = 12'hFFF;
            6629: color = 12'h888;
            6630: color = 12'h000;
            6631: color = 12'h000;
            6632: color = 12'h000;
            6633: color = 12'h000;
            6634: color = 12'h000;
            6635: color = 12'h000;
            6636: color = 12'h000;
            6637: color = 12'h000;
            6638: color = 12'h000;
            6639: color = 12'h000;
            6640: color = 12'h000;
            6641: color = 12'h888;
            6642: color = 12'hFFF;
            6643: color = 12'hFFF;
            6644: color = 12'hFFF;
            6645: color = 12'hFFF;
            6646: color = 12'hFFF;
            6647: color = 12'h777;
            6648: color = 12'h000;
            6649: color = 12'h000;
            6650: color = 12'h888;
            6651: color = 12'hFFF;
            6652: color = 12'hFFF;
            6653: color = 12'hFFF;
            6654: color = 12'hFFF;
            6655: color = 12'hFFF;
            6656: color = 12'hFFF;
            6657: color = 12'hFFF;
            6658: color = 12'hFFF;
            6659: color = 12'hFFF;
            6660: color = 12'hFFF;
            6661: color = 12'h000;
            6662: color = 12'h000;
            6663: color = 12'h000;
            6664: color = 12'h000;
            6665: color = 12'h888;
            6666: color = 12'hFFF;
            6667: color = 12'hFFF;
            6668: color = 12'h888;
            6669: color = 12'h111;
            6670: color = 12'hFFF;
            6671: color = 12'hFFF;
            6672: color = 12'hFFF;
            6673: color = 12'hFFF;
            6674: color = 12'h888;
            6675: color = 12'h000;
            6676: color = 12'h000;
            6677: color = 12'h888;
            6678: color = 12'hFFF;
            6679: color = 12'hFFF;
            6680: color = 12'hFFF;
            6681: color = 12'hFFF;
            6682: color = 12'hFFF;
            6683: color = 12'h777;
            6684: color = 12'h000;
            6685: color = 12'h000;
            6686: color = 12'h000;
            6687: color = 12'h000;
            6688: color = 12'h000;
            6689: color = 12'h000;
            6690: color = 12'h000;
            6691: color = 12'h000;
            6692: color = 12'h000;
            6693: color = 12'h000;
            6694: color = 12'h000;
            6695: color = 12'h000;
            6696: color = 12'h000;
            6697: color = 12'h000;
            6698: color = 12'h000;
            6699: color = 12'h000;
            6700: color = 12'h000;
            6701: color = 12'h000;
            6702: color = 12'h000;
            6703: color = 12'h000;
            6704: color = 12'h000;
            6705: color = 12'h000;
            6706: color = 12'h000;
            6707: color = 12'h000;
            6708: color = 12'h000;
            6709: color = 12'h000;
            6710: color = 12'h000;
            6711: color = 12'h000;
            6712: color = 12'h000;
            6713: color = 12'h000;
            6714: color = 12'h000;
            6715: color = 12'h000;
            6716: color = 12'h000;
            6717: color = 12'h000;
            6718: color = 12'h000;
            6719: color = 12'h000;
            6720: color = 12'h000;
            6721: color = 12'h000;
            6722: color = 12'h000;
            6723: color = 12'h000;
            6724: color = 12'h000;
            6725: color = 12'h000;
            6726: color = 12'h000;
            6727: color = 12'h000;
            6728: color = 12'h000;
            6729: color = 12'h000;
            6730: color = 12'h000;
            6731: color = 12'h000;
            6732: color = 12'h000;
            6733: color = 12'h000;
            6734: color = 12'h000;
            6735: color = 12'h000;
            6736: color = 12'h000;
            6737: color = 12'h000;
            6738: color = 12'h000;
            6739: color = 12'h000;
            6740: color = 12'h000;
            6741: color = 12'h000;
            6742: color = 12'h000;
            6743: color = 12'h000;
            6744: color = 12'h000;
            6745: color = 12'h000;
            6746: color = 12'h000;
            6747: color = 12'h000;
            6748: color = 12'h000;
            6749: color = 12'h000;
            6750: color = 12'h000;
            6751: color = 12'h000;
            6752: color = 12'h000;
            6753: color = 12'h000;
            6754: color = 12'h000;
            6755: color = 12'h000;
            6756: color = 12'h000;
            6757: color = 12'h000;
            6758: color = 12'h000;
            6759: color = 12'h000;
            6760: color = 12'h000;
            6761: color = 12'h000;
            6762: color = 12'h000;
            6763: color = 12'h000;
            6764: color = 12'h000;
            6765: color = 12'h000;
            6766: color = 12'h000;
            6767: color = 12'h000;
            6768: color = 12'h000;
            6769: color = 12'h888;
            6770: color = 12'hFFF;
            6771: color = 12'hFFF;
            6772: color = 12'hFFF;
            6773: color = 12'hFFF;
            6774: color = 12'hFFF;
            6775: color = 12'hFFF;
            6776: color = 12'hFFF;
            6777: color = 12'hFFF;
            6778: color = 12'hFFF;
            6779: color = 12'hFFF;
            6780: color = 12'hFFF;
            6781: color = 12'h888;
            6782: color = 12'h000;
            6783: color = 12'h000;
            6784: color = 12'h000;
            6785: color = 12'h000;
            6786: color = 12'hFFF;
            6787: color = 12'hFFF;
            6788: color = 12'hFFF;
            6789: color = 12'hFFF;
            6790: color = 12'hFFF;
            6791: color = 12'hFFF;
            6792: color = 12'hFFF;
            6793: color = 12'hFFF;
            6794: color = 12'hFFF;
            6795: color = 12'hFFF;
            6796: color = 12'h777;
            6797: color = 12'h000;
            6798: color = 12'h000;
            6799: color = 12'h000;
            6800: color = 12'h000;
            6801: color = 12'hFFF;
            6802: color = 12'hFFF;
            6803: color = 12'hFFF;
            6804: color = 12'hFFF;
            6805: color = 12'hFFF;
            6806: color = 12'hFFF;
            6807: color = 12'hFFF;
            6808: color = 12'hFFF;
            6809: color = 12'hFFF;
            6810: color = 12'h000;
            6811: color = 12'h777;
            6812: color = 12'hFFF;
            6813: color = 12'hFFF;
            6814: color = 12'h888;
            6815: color = 12'h000;
            6816: color = 12'h000;
            6817: color = 12'h000;
            6818: color = 12'h000;
            6819: color = 12'h000;
            6820: color = 12'h000;
            6821: color = 12'h000;
            6822: color = 12'h000;
            6823: color = 12'h777;
            6824: color = 12'hFFF;
            6825: color = 12'hFFF;
            6826: color = 12'h888;
            6827: color = 12'h000;
            6828: color = 12'h000;
            6829: color = 12'h000;
            6830: color = 12'h000;
            6831: color = 12'h000;
            6832: color = 12'h000;
            6833: color = 12'h000;
            6834: color = 12'h000;
            6835: color = 12'h000;
            6836: color = 12'h000;
            6837: color = 12'h000;
            6838: color = 12'h000;
            6839: color = 12'h000;
            6840: color = 12'h000;
            6841: color = 12'h000;
            6842: color = 12'h000;
            6843: color = 12'hFFF;
            6844: color = 12'hFFF;
            6845: color = 12'hFFF;
            6846: color = 12'hFFF;
            6847: color = 12'hFFF;
            6848: color = 12'hFFF;
            6849: color = 12'hFFF;
            6850: color = 12'h777;
            6851: color = 12'h000;
            6852: color = 12'h000;
            6853: color = 12'h000;
            6854: color = 12'h000;
            6855: color = 12'h000;
            6856: color = 12'h000;
            6857: color = 12'h000;
            6858: color = 12'h000;
            6859: color = 12'h888;
            6860: color = 12'hFFF;
            6861: color = 12'hFFF;
            6862: color = 12'hFFF;
            6863: color = 12'hFFF;
            6864: color = 12'hFFF;
            6865: color = 12'hFFF;
            6866: color = 12'hFFF;
            6867: color = 12'hFFF;
            6868: color = 12'hFFF;
            6869: color = 12'hFFF;
            6870: color = 12'h000;
            6871: color = 12'h000;
            6872: color = 12'h000;
            6873: color = 12'h000;
            6874: color = 12'h888;
            6875: color = 12'hFFF;
            6876: color = 12'hFFF;
            6877: color = 12'hFFF;
            6878: color = 12'hFFF;
            6879: color = 12'hFFF;
            6880: color = 12'h888;
            6881: color = 12'h000;
            6882: color = 12'h000;
            6883: color = 12'h000;
            6884: color = 12'h000;
            6885: color = 12'h000;
            6886: color = 12'h888;
            6887: color = 12'hFFF;
            6888: color = 12'hFFF;
            6889: color = 12'hFFF;
            6890: color = 12'hFFF;
            6891: color = 12'hFFF;
            6892: color = 12'hFFF;
            6893: color = 12'hFFF;
            6894: color = 12'hFFF;
            6895: color = 12'h777;
            6896: color = 12'h000;
            6897: color = 12'hFFF;
            6898: color = 12'hFFF;
            6899: color = 12'hFFF;
            6900: color = 12'hFFF;
            6901: color = 12'hFFF;
            6902: color = 12'hFFF;
            6903: color = 12'hFFF;
            6904: color = 12'hFFF;
            6905: color = 12'hFFF;
            6906: color = 12'hFFF;
            6907: color = 12'h777;
            6908: color = 12'h000;
            6909: color = 12'h000;
            6910: color = 12'h000;
            6911: color = 12'h000;
            6912: color = 12'h000;
            6913: color = 12'h000;
            6914: color = 12'h000;
            6915: color = 12'h000;
            6916: color = 12'h888;
            6917: color = 12'hFFF;
            6918: color = 12'hFFF;
            6919: color = 12'hFFF;
            6920: color = 12'hFFF;
            6921: color = 12'hFFF;
            6922: color = 12'h888;
            6923: color = 12'h000;
            6924: color = 12'h000;
            6925: color = 12'h000;
            6926: color = 12'h000;
            6927: color = 12'h000;
            6928: color = 12'h888;
            6929: color = 12'hFFF;
            6930: color = 12'hFFF;
            6931: color = 12'hFFF;
            6932: color = 12'hFFF;
            6933: color = 12'hFFF;
            6934: color = 12'h888;
            6935: color = 12'h000;
            6936: color = 12'h000;
            6937: color = 12'h000;
            6938: color = 12'h000;
            6939: color = 12'h000;
            6940: color = 12'h000;
            6941: color = 12'h000;
            6942: color = 12'h000;
            6943: color = 12'h000;
            6944: color = 12'h000;
            6945: color = 12'h000;
            6946: color = 12'h000;
            6947: color = 12'h000;
            6948: color = 12'h000;
            6949: color = 12'h888;
            6950: color = 12'hFFF;
            6951: color = 12'hFFF;
            6952: color = 12'hFFF;
            6953: color = 12'hFFF;
            6954: color = 12'hFFF;
            6955: color = 12'hFFF;
            6956: color = 12'hEEE;
            6957: color = 12'h000;
            6958: color = 12'h000;
            6959: color = 12'h000;
            6960: color = 12'h000;
            6961: color = 12'h888;
            6962: color = 12'hFFF;
            6963: color = 12'hFFF;
            6964: color = 12'hFFF;
            6965: color = 12'hFFF;
            6966: color = 12'hFFF;
            6967: color = 12'h888;
            6968: color = 12'h000;
            6969: color = 12'h000;
            6970: color = 12'h888;
            6971: color = 12'hFFF;
            6972: color = 12'hFFF;
            6973: color = 12'hFFF;
            6974: color = 12'hFFF;
            6975: color = 12'hFFF;
            6976: color = 12'hFFF;
            6977: color = 12'hFFF;
            6978: color = 12'hFFF;
            6979: color = 12'hFFF;
            6980: color = 12'hFFF;
            6981: color = 12'h000;
            6982: color = 12'h000;
            6983: color = 12'h000;
            6984: color = 12'h000;
            6985: color = 12'h888;
            6986: color = 12'hFFF;
            6987: color = 12'hFFF;
            6988: color = 12'hFFF;
            6989: color = 12'hFFF;
            6990: color = 12'hFFF;
            6991: color = 12'hFFF;
            6992: color = 12'hFFF;
            6993: color = 12'hFFF;
            6994: color = 12'hFFF;
            6995: color = 12'hEEE;
            6996: color = 12'h000;
            6997: color = 12'h888;
            6998: color = 12'hFFF;
            6999: color = 12'hFFF;
            7000: color = 12'hFFF;
            7001: color = 12'hFFF;
            7002: color = 12'hFFF;
            7003: color = 12'h888;
            7004: color = 12'h000;
            7005: color = 12'h000;
            7006: color = 12'h000;
            7007: color = 12'h000;
            7008: color = 12'h000;
            7009: color = 12'h000;
            7010: color = 12'h000;
            7011: color = 12'h000;
            7012: color = 12'h000;
            7013: color = 12'h000;
            7014: color = 12'h000;
            7015: color = 12'h000;
            7016: color = 12'h000;
            7017: color = 12'h000;
            7018: color = 12'h000;
            7019: color = 12'h000;
            7020: color = 12'h000;
            7021: color = 12'h000;
            7022: color = 12'h000;
            7023: color = 12'h000;
            7024: color = 12'h000;
            7025: color = 12'h000;
            7026: color = 12'h000;
            7027: color = 12'h000;
            7028: color = 12'h000;
            7029: color = 12'h000;
            7030: color = 12'h000;
            7031: color = 12'h000;
            7032: color = 12'h000;
            7033: color = 12'h000;
            7034: color = 12'h000;
            7035: color = 12'h000;
            7036: color = 12'h000;
            7037: color = 12'h000;
            7038: color = 12'h000;
            7039: color = 12'h000;
            7040: color = 12'h000;
            7041: color = 12'h000;
            7042: color = 12'h000;
            7043: color = 12'h000;
            7044: color = 12'h000;
            7045: color = 12'h000;
            7046: color = 12'h000;
            7047: color = 12'h000;
            7048: color = 12'h000;
            7049: color = 12'h000;
            7050: color = 12'h000;
            7051: color = 12'h000;
            7052: color = 12'h000;
            7053: color = 12'h000;
            7054: color = 12'h000;
            7055: color = 12'h000;
            7056: color = 12'h000;
            7057: color = 12'h000;
            7058: color = 12'h000;
            7059: color = 12'h000;
            7060: color = 12'h000;
            7061: color = 12'h000;
            7062: color = 12'h000;
            7063: color = 12'h000;
            7064: color = 12'h000;
            7065: color = 12'h000;
            7066: color = 12'h000;
            7067: color = 12'h000;
            7068: color = 12'h000;
            7069: color = 12'h000;
            7070: color = 12'h000;
            7071: color = 12'h000;
            7072: color = 12'h000;
            7073: color = 12'h000;
            7074: color = 12'h000;
            7075: color = 12'h000;
            7076: color = 12'h000;
            7077: color = 12'h000;
            7078: color = 12'h000;
            7079: color = 12'h000;
            7080: color = 12'h000;
            7081: color = 12'h000;
            7082: color = 12'h000;
            7083: color = 12'h000;
            7084: color = 12'h000;
            7085: color = 12'h000;
            7086: color = 12'h000;
            7087: color = 12'h000;
            7088: color = 12'h000;
            7089: color = 12'h888;
            7090: color = 12'hFFF;
            7091: color = 12'hFFF;
            7092: color = 12'hFFF;
            7093: color = 12'hFFF;
            7094: color = 12'hFFF;
            7095: color = 12'hFFF;
            7096: color = 12'hFFF;
            7097: color = 12'hFFF;
            7098: color = 12'hFFF;
            7099: color = 12'hFFF;
            7100: color = 12'hFFF;
            7101: color = 12'h777;
            7102: color = 12'h000;
            7103: color = 12'h000;
            7104: color = 12'h000;
            7105: color = 12'h000;
            7106: color = 12'hFFF;
            7107: color = 12'hFFF;
            7108: color = 12'hFFF;
            7109: color = 12'hFFF;
            7110: color = 12'hCCC;
            7111: color = 12'h888;
            7112: color = 12'h888;
            7113: color = 12'h888;
            7114: color = 12'h888;
            7115: color = 12'hFFF;
            7116: color = 12'h777;
            7117: color = 12'h000;
            7118: color = 12'h777;
            7119: color = 12'h888;
            7120: color = 12'h888;
            7121: color = 12'h888;
            7122: color = 12'h888;
            7123: color = 12'h888;
            7124: color = 12'h888;
            7125: color = 12'h888;
            7126: color = 12'h888;
            7127: color = 12'hFFF;
            7128: color = 12'hFFF;
            7129: color = 12'hFFF;
            7130: color = 12'h000;
            7131: color = 12'h888;
            7132: color = 12'hFFF;
            7133: color = 12'hFFF;
            7134: color = 12'h777;
            7135: color = 12'h000;
            7136: color = 12'h000;
            7137: color = 12'h000;
            7138: color = 12'h000;
            7139: color = 12'h000;
            7140: color = 12'h000;
            7141: color = 12'h000;
            7142: color = 12'h000;
            7143: color = 12'h888;
            7144: color = 12'hFFF;
            7145: color = 12'hFFF;
            7146: color = 12'h777;
            7147: color = 12'h000;
            7148: color = 12'h000;
            7149: color = 12'h000;
            7150: color = 12'h000;
            7151: color = 12'h000;
            7152: color = 12'h000;
            7153: color = 12'h000;
            7154: color = 12'h000;
            7155: color = 12'h000;
            7156: color = 12'h000;
            7157: color = 12'h000;
            7158: color = 12'h000;
            7159: color = 12'h000;
            7160: color = 12'h000;
            7161: color = 12'h000;
            7162: color = 12'h000;
            7163: color = 12'hFFF;
            7164: color = 12'hFFF;
            7165: color = 12'hFFF;
            7166: color = 12'hFFF;
            7167: color = 12'hFFF;
            7168: color = 12'hFFF;
            7169: color = 12'hFFF;
            7170: color = 12'h777;
            7171: color = 12'h000;
            7172: color = 12'h000;
            7173: color = 12'h000;
            7174: color = 12'h000;
            7175: color = 12'h000;
            7176: color = 12'h000;
            7177: color = 12'h000;
            7178: color = 12'h000;
            7179: color = 12'h888;
            7180: color = 12'hFFF;
            7181: color = 12'hFFF;
            7182: color = 12'hCCC;
            7183: color = 12'h888;
            7184: color = 12'h888;
            7185: color = 12'h888;
            7186: color = 12'h888;
            7187: color = 12'h888;
            7188: color = 12'h888;
            7189: color = 12'h888;
            7190: color = 12'h888;
            7191: color = 12'h888;
            7192: color = 12'h777;
            7193: color = 12'h000;
            7194: color = 12'h444;
            7195: color = 12'h888;
            7196: color = 12'hFFF;
            7197: color = 12'hFFF;
            7198: color = 12'hFFF;
            7199: color = 12'h888;
            7200: color = 12'h444;
            7201: color = 12'h000;
            7202: color = 12'h000;
            7203: color = 12'h444;
            7204: color = 12'h888;
            7205: color = 12'h888;
            7206: color = 12'h888;
            7207: color = 12'h888;
            7208: color = 12'h888;
            7209: color = 12'h888;
            7210: color = 12'h888;
            7211: color = 12'h888;
            7212: color = 12'hCCC;
            7213: color = 12'hFFF;
            7214: color = 12'hFFF;
            7215: color = 12'h777;
            7216: color = 12'h000;
            7217: color = 12'hFFF;
            7218: color = 12'hFFF;
            7219: color = 12'hFFF;
            7220: color = 12'hFFF;
            7221: color = 12'hCCC;
            7222: color = 12'h888;
            7223: color = 12'h888;
            7224: color = 12'h888;
            7225: color = 12'h888;
            7226: color = 12'hFFF;
            7227: color = 12'h777;
            7228: color = 12'h000;
            7229: color = 12'h000;
            7230: color = 12'h000;
            7231: color = 12'h000;
            7232: color = 12'h000;
            7233: color = 12'h000;
            7234: color = 12'h000;
            7235: color = 12'h000;
            7236: color = 12'h444;
            7237: color = 12'h888;
            7238: color = 12'hFFF;
            7239: color = 12'hFFF;
            7240: color = 12'hFFF;
            7241: color = 12'h888;
            7242: color = 12'h444;
            7243: color = 12'h000;
            7244: color = 12'h000;
            7245: color = 12'h444;
            7246: color = 12'h888;
            7247: color = 12'h888;
            7248: color = 12'h888;
            7249: color = 12'h888;
            7250: color = 12'h888;
            7251: color = 12'h888;
            7252: color = 12'h888;
            7253: color = 12'h888;
            7254: color = 12'h888;
            7255: color = 12'h888;
            7256: color = 12'h888;
            7257: color = 12'h444;
            7258: color = 12'h000;
            7259: color = 12'h000;
            7260: color = 12'h000;
            7261: color = 12'h000;
            7262: color = 12'h000;
            7263: color = 12'h000;
            7264: color = 12'h000;
            7265: color = 12'h000;
            7266: color = 12'h000;
            7267: color = 12'h000;
            7268: color = 12'h000;
            7269: color = 12'h888;
            7270: color = 12'hFFF;
            7271: color = 12'hFFF;
            7272: color = 12'hFFF;
            7273: color = 12'hFFF;
            7274: color = 12'hFFF;
            7275: color = 12'hFFF;
            7276: color = 12'hFFF;
            7277: color = 12'h000;
            7278: color = 12'h000;
            7279: color = 12'h000;
            7280: color = 12'h000;
            7281: color = 12'h444;
            7282: color = 12'h888;
            7283: color = 12'hFFF;
            7284: color = 12'hFFF;
            7285: color = 12'hFFF;
            7286: color = 12'h888;
            7287: color = 12'h444;
            7288: color = 12'h000;
            7289: color = 12'h000;
            7290: color = 12'h444;
            7291: color = 12'h888;
            7292: color = 12'h888;
            7293: color = 12'h888;
            7294: color = 12'h888;
            7295: color = 12'h888;
            7296: color = 12'h888;
            7297: color = 12'h888;
            7298: color = 12'h888;
            7299: color = 12'h888;
            7300: color = 12'h888;
            7301: color = 12'h888;
            7302: color = 12'h888;
            7303: color = 12'h777;
            7304: color = 12'h000;
            7305: color = 12'h888;
            7306: color = 12'hFFF;
            7307: color = 12'hFFF;
            7308: color = 12'hFFF;
            7309: color = 12'hFFF;
            7310: color = 12'h888;
            7311: color = 12'h888;
            7312: color = 12'h888;
            7313: color = 12'h888;
            7314: color = 12'hCCC;
            7315: color = 12'hFFF;
            7316: color = 12'h000;
            7317: color = 12'h444;
            7318: color = 12'h888;
            7319: color = 12'hFFF;
            7320: color = 12'hFFF;
            7321: color = 12'hFFF;
            7322: color = 12'h888;
            7323: color = 12'h444;
            7324: color = 12'h000;
            7325: color = 12'h000;
            7326: color = 12'h000;
            7327: color = 12'h000;
            7328: color = 12'h000;
            7329: color = 12'h000;
            7330: color = 12'h000;
            7331: color = 12'h000;
            7332: color = 12'h000;
            7333: color = 12'h000;
            7334: color = 12'h000;
            7335: color = 12'h000;
            7336: color = 12'h000;
            7337: color = 12'h000;
            7338: color = 12'h000;
            7339: color = 12'h000;
            7340: color = 12'h000;
            7341: color = 12'h000;
            7342: color = 12'h000;
            7343: color = 12'h000;
            7344: color = 12'h000;
            7345: color = 12'h000;
            7346: color = 12'h000;
            7347: color = 12'h000;
            7348: color = 12'h000;
            7349: color = 12'h000;
            7350: color = 12'h000;
            7351: color = 12'h000;
            7352: color = 12'h000;
            7353: color = 12'h000;
            7354: color = 12'h000;
            7355: color = 12'h000;
            7356: color = 12'h000;
            7357: color = 12'h000;
            7358: color = 12'h000;
            7359: color = 12'h000;
            7360: color = 12'h000;
            7361: color = 12'h000;
            7362: color = 12'h000;
            7363: color = 12'h000;
            7364: color = 12'h000;
            7365: color = 12'h000;
            7366: color = 12'h000;
            7367: color = 12'h000;
            7368: color = 12'h000;
            7369: color = 12'h000;
            7370: color = 12'h000;
            7371: color = 12'h000;
            7372: color = 12'h000;
            7373: color = 12'h000;
            7374: color = 12'h000;
            7375: color = 12'h000;
            7376: color = 12'h000;
            7377: color = 12'h000;
            7378: color = 12'h000;
            7379: color = 12'h000;
            7380: color = 12'h000;
            7381: color = 12'h000;
            7382: color = 12'h000;
            7383: color = 12'h000;
            7384: color = 12'h000;
            7385: color = 12'h000;
            7386: color = 12'h000;
            7387: color = 12'h000;
            7388: color = 12'h000;
            7389: color = 12'h000;
            7390: color = 12'h000;
            7391: color = 12'h000;
            7392: color = 12'h000;
            7393: color = 12'h000;
            7394: color = 12'h000;
            7395: color = 12'h000;
            7396: color = 12'h000;
            7397: color = 12'h000;
            7398: color = 12'h000;
            7399: color = 12'h000;
            7400: color = 12'h000;
            7401: color = 12'h000;
            7402: color = 12'h000;
            7403: color = 12'h000;
            7404: color = 12'h000;
            7405: color = 12'h000;
            7406: color = 12'h000;
            7407: color = 12'h000;
            7408: color = 12'h000;
            7409: color = 12'h888;
            7410: color = 12'hFFF;
            7411: color = 12'hFFF;
            7412: color = 12'hFFF;
            7413: color = 12'hFFF;
            7414: color = 12'hFFF;
            7415: color = 12'hFFF;
            7416: color = 12'hFFF;
            7417: color = 12'hFFF;
            7418: color = 12'hFFF;
            7419: color = 12'hFFF;
            7420: color = 12'hFFF;
            7421: color = 12'h777;
            7422: color = 12'h000;
            7423: color = 12'h000;
            7424: color = 12'h000;
            7425: color = 12'h000;
            7426: color = 12'hFFF;
            7427: color = 12'hFFF;
            7428: color = 12'hFFF;
            7429: color = 12'hFFF;
            7430: color = 12'h777;
            7431: color = 12'h000;
            7432: color = 12'h000;
            7433: color = 12'h000;
            7434: color = 12'h000;
            7435: color = 12'hEEE;
            7436: color = 12'h777;
            7437: color = 12'h000;
            7438: color = 12'hFFF;
            7439: color = 12'hFFF;
            7440: color = 12'hFFF;
            7441: color = 12'h111;
            7442: color = 12'h000;
            7443: color = 12'h000;
            7444: color = 12'h000;
            7445: color = 12'h000;
            7446: color = 12'h111;
            7447: color = 12'hFFF;
            7448: color = 12'hFFF;
            7449: color = 12'hFFF;
            7450: color = 12'h000;
            7451: color = 12'h777;
            7452: color = 12'hFFF;
            7453: color = 12'hFFF;
            7454: color = 12'h888;
            7455: color = 12'h000;
            7456: color = 12'h000;
            7457: color = 12'h000;
            7458: color = 12'h000;
            7459: color = 12'h000;
            7460: color = 12'h000;
            7461: color = 12'h000;
            7462: color = 12'h000;
            7463: color = 12'h777;
            7464: color = 12'hFFF;
            7465: color = 12'hFFF;
            7466: color = 12'h888;
            7467: color = 12'h000;
            7468: color = 12'h000;
            7469: color = 12'h000;
            7470: color = 12'h000;
            7471: color = 12'h000;
            7472: color = 12'h000;
            7473: color = 12'h000;
            7474: color = 12'h000;
            7475: color = 12'h000;
            7476: color = 12'h000;
            7477: color = 12'h000;
            7478: color = 12'h000;
            7479: color = 12'h000;
            7480: color = 12'h000;
            7481: color = 12'h000;
            7482: color = 12'h000;
            7483: color = 12'hFFF;
            7484: color = 12'hFFF;
            7485: color = 12'hFFF;
            7486: color = 12'hFFF;
            7487: color = 12'hFFF;
            7488: color = 12'hFFF;
            7489: color = 12'hFFF;
            7490: color = 12'h777;
            7491: color = 12'h000;
            7492: color = 12'h000;
            7493: color = 12'h000;
            7494: color = 12'h000;
            7495: color = 12'h000;
            7496: color = 12'h000;
            7497: color = 12'h000;
            7498: color = 12'h000;
            7499: color = 12'h888;
            7500: color = 12'hFFF;
            7501: color = 12'hFFF;
            7502: color = 12'h777;
            7503: color = 12'h000;
            7504: color = 12'h000;
            7505: color = 12'h000;
            7506: color = 12'h000;
            7507: color = 12'h000;
            7508: color = 12'h000;
            7509: color = 12'h000;
            7510: color = 12'hFFF;
            7511: color = 12'hFFF;
            7512: color = 12'hFFF;
            7513: color = 12'h000;
            7514: color = 12'h000;
            7515: color = 12'h000;
            7516: color = 12'hFFF;
            7517: color = 12'hFFF;
            7518: color = 12'hFFF;
            7519: color = 12'h000;
            7520: color = 12'h000;
            7521: color = 12'h000;
            7522: color = 12'h000;
            7523: color = 12'h888;
            7524: color = 12'hFFF;
            7525: color = 12'hFFF;
            7526: color = 12'h888;
            7527: color = 12'h000;
            7528: color = 12'h000;
            7529: color = 12'h000;
            7530: color = 12'h000;
            7531: color = 12'h000;
            7532: color = 12'h888;
            7533: color = 12'hFFF;
            7534: color = 12'hFFF;
            7535: color = 12'h777;
            7536: color = 12'h000;
            7537: color = 12'hFFF;
            7538: color = 12'hFFF;
            7539: color = 12'hFFF;
            7540: color = 12'hFFF;
            7541: color = 12'h777;
            7542: color = 12'h000;
            7543: color = 12'h000;
            7544: color = 12'h000;
            7545: color = 12'h000;
            7546: color = 12'hEEE;
            7547: color = 12'h777;
            7548: color = 12'h000;
            7549: color = 12'h000;
            7550: color = 12'h000;
            7551: color = 12'h000;
            7552: color = 12'h000;
            7553: color = 12'h000;
            7554: color = 12'h000;
            7555: color = 12'h000;
            7556: color = 12'h000;
            7557: color = 12'h000;
            7558: color = 12'hFFF;
            7559: color = 12'hFFF;
            7560: color = 12'hFFF;
            7561: color = 12'h000;
            7562: color = 12'h000;
            7563: color = 12'h000;
            7564: color = 12'h000;
            7565: color = 12'h888;
            7566: color = 12'hFFF;
            7567: color = 12'hFFF;
            7568: color = 12'h777;
            7569: color = 12'h000;
            7570: color = 12'h000;
            7571: color = 12'h000;
            7572: color = 12'h000;
            7573: color = 12'h000;
            7574: color = 12'h888;
            7575: color = 12'hFFF;
            7576: color = 12'hFFF;
            7577: color = 12'h777;
            7578: color = 12'h000;
            7579: color = 12'h000;
            7580: color = 12'h000;
            7581: color = 12'h000;
            7582: color = 12'h000;
            7583: color = 12'h000;
            7584: color = 12'h000;
            7585: color = 12'h000;
            7586: color = 12'h000;
            7587: color = 12'h000;
            7588: color = 12'h000;
            7589: color = 12'h777;
            7590: color = 12'hFFF;
            7591: color = 12'hFFF;
            7592: color = 12'hFFF;
            7593: color = 12'hFFF;
            7594: color = 12'hFFF;
            7595: color = 12'hFFF;
            7596: color = 12'hEEE;
            7597: color = 12'h111;
            7598: color = 12'h000;
            7599: color = 12'h000;
            7600: color = 12'h000;
            7601: color = 12'h000;
            7602: color = 12'h000;
            7603: color = 12'hFFF;
            7604: color = 12'hFFF;
            7605: color = 12'hFFF;
            7606: color = 12'h000;
            7607: color = 12'h000;
            7608: color = 12'h000;
            7609: color = 12'h000;
            7610: color = 12'h000;
            7611: color = 12'h000;
            7612: color = 12'h000;
            7613: color = 12'h000;
            7614: color = 12'h000;
            7615: color = 12'h000;
            7616: color = 12'h000;
            7617: color = 12'h000;
            7618: color = 12'h000;
            7619: color = 12'h000;
            7620: color = 12'h111;
            7621: color = 12'hFFF;
            7622: color = 12'hFFF;
            7623: color = 12'hFFF;
            7624: color = 12'h000;
            7625: color = 12'h888;
            7626: color = 12'hFFF;
            7627: color = 12'hFFF;
            7628: color = 12'hFFF;
            7629: color = 12'hEEE;
            7630: color = 12'h000;
            7631: color = 12'h000;
            7632: color = 12'h000;
            7633: color = 12'h000;
            7634: color = 12'h888;
            7635: color = 12'hEEE;
            7636: color = 12'h000;
            7637: color = 12'h000;
            7638: color = 12'h000;
            7639: color = 12'hFFF;
            7640: color = 12'hFFF;
            7641: color = 12'hFFF;
            7642: color = 12'h000;
            7643: color = 12'h000;
            7644: color = 12'h000;
            7645: color = 12'h000;
            7646: color = 12'h000;
            7647: color = 12'h000;
            7648: color = 12'h000;
            7649: color = 12'h000;
            7650: color = 12'h000;
            7651: color = 12'h000;
            7652: color = 12'h000;
            7653: color = 12'h000;
            7654: color = 12'h000;
            7655: color = 12'h000;
            7656: color = 12'h000;
            7657: color = 12'h000;
            7658: color = 12'h000;
            7659: color = 12'h000;
            7660: color = 12'h000;
            7661: color = 12'h000;
            7662: color = 12'h000;
            7663: color = 12'h000;
            7664: color = 12'h000;
            7665: color = 12'h000;
            7666: color = 12'h000;
            7667: color = 12'h000;
            7668: color = 12'h000;
            7669: color = 12'h000;
            7670: color = 12'h000;
            7671: color = 12'h000;
            7672: color = 12'h000;
            7673: color = 12'h000;
            7674: color = 12'h000;
            7675: color = 12'h000;
            7676: color = 12'h000;
            7677: color = 12'h000;
            7678: color = 12'h000;
            7679: color = 12'h000;
            7680: color = 12'h000;
            7681: color = 12'h000;
            7682: color = 12'h000;
            7683: color = 12'h000;
            7684: color = 12'h000;
            7685: color = 12'h000;
            7686: color = 12'h000;
            7687: color = 12'h000;
            7688: color = 12'h000;
            7689: color = 12'h000;
            7690: color = 12'h000;
            7691: color = 12'h000;
            7692: color = 12'h000;
            7693: color = 12'h000;
            7694: color = 12'h000;
            7695: color = 12'h000;
            7696: color = 12'h000;
            7697: color = 12'h000;
            7698: color = 12'h000;
            7699: color = 12'h000;
            7700: color = 12'h000;
            7701: color = 12'h000;
            7702: color = 12'h000;
            7703: color = 12'h000;
            7704: color = 12'h000;
            7705: color = 12'h000;
            7706: color = 12'h000;
            7707: color = 12'h000;
            7708: color = 12'h000;
            7709: color = 12'h000;
            7710: color = 12'h000;
            7711: color = 12'h000;
            7712: color = 12'h000;
            7713: color = 12'h000;
            7714: color = 12'h000;
            7715: color = 12'h000;
            7716: color = 12'h000;
            7717: color = 12'h000;
            7718: color = 12'h000;
            7719: color = 12'h000;
            7720: color = 12'h000;
            7721: color = 12'h000;
            7722: color = 12'h000;
            7723: color = 12'h000;
            7724: color = 12'h000;
            7725: color = 12'h000;
            7726: color = 12'h000;
            7727: color = 12'h000;
            7728: color = 12'h000;
            7729: color = 12'h888;
            7730: color = 12'hFFF;
            7731: color = 12'hFFF;
            7732: color = 12'h888;
            7733: color = 12'h000;
            7734: color = 12'h000;
            7735: color = 12'h000;
            7736: color = 12'h000;
            7737: color = 12'h000;
            7738: color = 12'h000;
            7739: color = 12'h000;
            7740: color = 12'h000;
            7741: color = 12'h000;
            7742: color = 12'h000;
            7743: color = 12'h000;
            7744: color = 12'h000;
            7745: color = 12'h000;
            7746: color = 12'hFFF;
            7747: color = 12'hFFF;
            7748: color = 12'hFFF;
            7749: color = 12'h111;
            7750: color = 12'h000;
            7751: color = 12'h000;
            7752: color = 12'h000;
            7753: color = 12'h000;
            7754: color = 12'h000;
            7755: color = 12'h000;
            7756: color = 12'h000;
            7757: color = 12'h000;
            7758: color = 12'hFFF;
            7759: color = 12'hFFF;
            7760: color = 12'hFFF;
            7761: color = 12'hFFF;
            7762: color = 12'hFFF;
            7763: color = 12'hFFF;
            7764: color = 12'hFFF;
            7765: color = 12'hFFF;
            7766: color = 12'hFFF;
            7767: color = 12'hFFF;
            7768: color = 12'hFFF;
            7769: color = 12'hFFF;
            7770: color = 12'h000;
            7771: color = 12'h000;
            7772: color = 12'h000;
            7773: color = 12'h000;
            7774: color = 12'h888;
            7775: color = 12'hFFF;
            7776: color = 12'hFFF;
            7777: color = 12'hFFF;
            7778: color = 12'hEEE;
            7779: color = 12'h000;
            7780: color = 12'h000;
            7781: color = 12'h000;
            7782: color = 12'h000;
            7783: color = 12'h000;
            7784: color = 12'h000;
            7785: color = 12'h000;
            7786: color = 12'h888;
            7787: color = 12'hFFF;
            7788: color = 12'hFFF;
            7789: color = 12'hFFF;
            7790: color = 12'hEEE;
            7791: color = 12'h000;
            7792: color = 12'h000;
            7793: color = 12'h000;
            7794: color = 12'h000;
            7795: color = 12'h000;
            7796: color = 12'h000;
            7797: color = 12'h000;
            7798: color = 12'h000;
            7799: color = 12'h000;
            7800: color = 12'h000;
            7801: color = 12'h000;
            7802: color = 12'h000;
            7803: color = 12'hFFF;
            7804: color = 12'hFFF;
            7805: color = 12'hFFF;
            7806: color = 12'h111;
            7807: color = 12'h000;
            7808: color = 12'h000;
            7809: color = 12'h000;
            7810: color = 12'h000;
            7811: color = 12'h000;
            7812: color = 12'h000;
            7813: color = 12'h000;
            7814: color = 12'h000;
            7815: color = 12'h000;
            7816: color = 12'h000;
            7817: color = 12'h000;
            7818: color = 12'h000;
            7819: color = 12'h888;
            7820: color = 12'hFFF;
            7821: color = 12'hFFF;
            7822: color = 12'h777;
            7823: color = 12'h000;
            7824: color = 12'h000;
            7825: color = 12'h000;
            7826: color = 12'h000;
            7827: color = 12'h000;
            7828: color = 12'h000;
            7829: color = 12'h000;
            7830: color = 12'hFFF;
            7831: color = 12'hFFF;
            7832: color = 12'hFFF;
            7833: color = 12'h000;
            7834: color = 12'h000;
            7835: color = 12'h000;
            7836: color = 12'hFFF;
            7837: color = 12'hFFF;
            7838: color = 12'hFFF;
            7839: color = 12'h000;
            7840: color = 12'h000;
            7841: color = 12'h000;
            7842: color = 12'h000;
            7843: color = 12'h888;
            7844: color = 12'hFFF;
            7845: color = 12'hFFF;
            7846: color = 12'hFFF;
            7847: color = 12'hFFF;
            7848: color = 12'hFFF;
            7849: color = 12'hFFF;
            7850: color = 12'hFFF;
            7851: color = 12'hFFF;
            7852: color = 12'hFFF;
            7853: color = 12'hFFF;
            7854: color = 12'hFFF;
            7855: color = 12'h888;
            7856: color = 12'h000;
            7857: color = 12'hFFF;
            7858: color = 12'hFFF;
            7859: color = 12'hFFF;
            7860: color = 12'h111;
            7861: color = 12'h000;
            7862: color = 12'h000;
            7863: color = 12'h000;
            7864: color = 12'h000;
            7865: color = 12'h000;
            7866: color = 12'h000;
            7867: color = 12'h000;
            7868: color = 12'h000;
            7869: color = 12'h000;
            7870: color = 12'h000;
            7871: color = 12'h000;
            7872: color = 12'h000;
            7873: color = 12'h000;
            7874: color = 12'h000;
            7875: color = 12'h000;
            7876: color = 12'h000;
            7877: color = 12'h000;
            7878: color = 12'hFFF;
            7879: color = 12'hFFF;
            7880: color = 12'hFFF;
            7881: color = 12'h000;
            7882: color = 12'h000;
            7883: color = 12'h000;
            7884: color = 12'h000;
            7885: color = 12'h888;
            7886: color = 12'hFFF;
            7887: color = 12'hFFF;
            7888: color = 12'h777;
            7889: color = 12'h000;
            7890: color = 12'h000;
            7891: color = 12'h000;
            7892: color = 12'h000;
            7893: color = 12'h000;
            7894: color = 12'h888;
            7895: color = 12'hFFF;
            7896: color = 12'hFFF;
            7897: color = 12'h777;
            7898: color = 12'h000;
            7899: color = 12'h000;
            7900: color = 12'h000;
            7901: color = 12'h000;
            7902: color = 12'h000;
            7903: color = 12'h000;
            7904: color = 12'h000;
            7905: color = 12'h000;
            7906: color = 12'h000;
            7907: color = 12'h000;
            7908: color = 12'h000;
            7909: color = 12'h000;
            7910: color = 12'h000;
            7911: color = 12'h000;
            7912: color = 12'h000;
            7913: color = 12'h000;
            7914: color = 12'h000;
            7915: color = 12'h000;
            7916: color = 12'h111;
            7917: color = 12'hEEE;
            7918: color = 12'hFFF;
            7919: color = 12'hEEE;
            7920: color = 12'h000;
            7921: color = 12'h000;
            7922: color = 12'h000;
            7923: color = 12'hFFF;
            7924: color = 12'hFFF;
            7925: color = 12'hFFF;
            7926: color = 12'h000;
            7927: color = 12'h000;
            7928: color = 12'h000;
            7929: color = 12'h000;
            7930: color = 12'h000;
            7931: color = 12'h000;
            7932: color = 12'h000;
            7933: color = 12'h777;
            7934: color = 12'hFFF;
            7935: color = 12'hFFF;
            7936: color = 12'hFFF;
            7937: color = 12'hFFF;
            7938: color = 12'hFFF;
            7939: color = 12'hFFF;
            7940: color = 12'hFFF;
            7941: color = 12'hFFF;
            7942: color = 12'hFFF;
            7943: color = 12'hFFF;
            7944: color = 12'h000;
            7945: color = 12'h888;
            7946: color = 12'hFFF;
            7947: color = 12'hFFF;
            7948: color = 12'h888;
            7949: color = 12'h000;
            7950: color = 12'h000;
            7951: color = 12'h000;
            7952: color = 12'h000;
            7953: color = 12'h000;
            7954: color = 12'h000;
            7955: color = 12'h000;
            7956: color = 12'h000;
            7957: color = 12'h000;
            7958: color = 12'h000;
            7959: color = 12'hFFF;
            7960: color = 12'hFFF;
            7961: color = 12'hFFF;
            7962: color = 12'h000;
            7963: color = 12'h000;
            7964: color = 12'h000;
            7965: color = 12'h000;
            7966: color = 12'h000;
            7967: color = 12'h000;
            7968: color = 12'h000;
            7969: color = 12'h000;
            7970: color = 12'h000;
            7971: color = 12'h000;
            7972: color = 12'h000;
            7973: color = 12'h000;
            7974: color = 12'h000;
            7975: color = 12'h000;
            7976: color = 12'h000;
            7977: color = 12'h000;
            7978: color = 12'h000;
            7979: color = 12'h000;
            7980: color = 12'h000;
            7981: color = 12'h000;
            7982: color = 12'h000;
            7983: color = 12'h000;
            7984: color = 12'h000;
            7985: color = 12'h000;
            7986: color = 12'h000;
            7987: color = 12'h000;
            7988: color = 12'h000;
            7989: color = 12'h000;
            7990: color = 12'h000;
            7991: color = 12'h000;
            7992: color = 12'h000;
            7993: color = 12'h000;
            7994: color = 12'h000;
            7995: color = 12'h000;
            7996: color = 12'h000;
            7997: color = 12'h000;
            7998: color = 12'h000;
            7999: color = 12'h000;
            8000: color = 12'h000;
            8001: color = 12'h000;
            8002: color = 12'h000;
            8003: color = 12'h000;
            8004: color = 12'h000;
            8005: color = 12'h000;
            8006: color = 12'h000;
            8007: color = 12'h000;
            8008: color = 12'h000;
            8009: color = 12'h000;
            8010: color = 12'h000;
            8011: color = 12'h000;
            8012: color = 12'h000;
            8013: color = 12'h000;
            8014: color = 12'h000;
            8015: color = 12'h000;
            8016: color = 12'h000;
            8017: color = 12'h000;
            8018: color = 12'h000;
            8019: color = 12'h000;
            8020: color = 12'h000;
            8021: color = 12'h000;
            8022: color = 12'h000;
            8023: color = 12'h000;
            8024: color = 12'h000;
            8025: color = 12'h000;
            8026: color = 12'h000;
            8027: color = 12'h000;
            8028: color = 12'h000;
            8029: color = 12'h000;
            8030: color = 12'h000;
            8031: color = 12'h000;
            8032: color = 12'h000;
            8033: color = 12'h000;
            8034: color = 12'h000;
            8035: color = 12'h000;
            8036: color = 12'h000;
            8037: color = 12'h000;
            8038: color = 12'h000;
            8039: color = 12'h000;
            8040: color = 12'h000;
            8041: color = 12'h000;
            8042: color = 12'h000;
            8043: color = 12'h000;
            8044: color = 12'h000;
            8045: color = 12'h000;
            8046: color = 12'h000;
            8047: color = 12'h000;
            8048: color = 12'h000;
            8049: color = 12'h888;
            8050: color = 12'hFFF;
            8051: color = 12'hFFF;
            8052: color = 12'h777;
            8053: color = 12'h000;
            8054: color = 12'h000;
            8055: color = 12'h000;
            8056: color = 12'h000;
            8057: color = 12'h000;
            8058: color = 12'h000;
            8059: color = 12'h000;
            8060: color = 12'h000;
            8061: color = 12'h000;
            8062: color = 12'h000;
            8063: color = 12'h000;
            8064: color = 12'h000;
            8065: color = 12'h000;
            8066: color = 12'hFFF;
            8067: color = 12'hFFF;
            8068: color = 12'hFFF;
            8069: color = 12'h000;
            8070: color = 12'h000;
            8071: color = 12'h000;
            8072: color = 12'h000;
            8073: color = 12'h000;
            8074: color = 12'h000;
            8075: color = 12'h000;
            8076: color = 12'h000;
            8077: color = 12'h000;
            8078: color = 12'hFFF;
            8079: color = 12'hFFF;
            8080: color = 12'hFFF;
            8081: color = 12'hFFF;
            8082: color = 12'hFFF;
            8083: color = 12'hFFF;
            8084: color = 12'hFFF;
            8085: color = 12'hFFF;
            8086: color = 12'hFFF;
            8087: color = 12'h888;
            8088: color = 12'h888;
            8089: color = 12'h777;
            8090: color = 12'h000;
            8091: color = 12'h000;
            8092: color = 12'h000;
            8093: color = 12'h000;
            8094: color = 12'h888;
            8095: color = 12'hFFF;
            8096: color = 12'hFFF;
            8097: color = 12'hFFF;
            8098: color = 12'hFFF;
            8099: color = 12'h000;
            8100: color = 12'h000;
            8101: color = 12'h000;
            8102: color = 12'h000;
            8103: color = 12'h000;
            8104: color = 12'h000;
            8105: color = 12'h000;
            8106: color = 12'h888;
            8107: color = 12'hFFF;
            8108: color = 12'hFFF;
            8109: color = 12'hFFF;
            8110: color = 12'hFFF;
            8111: color = 12'h000;
            8112: color = 12'h000;
            8113: color = 12'h000;
            8114: color = 12'h000;
            8115: color = 12'h000;
            8116: color = 12'h000;
            8117: color = 12'h000;
            8118: color = 12'h000;
            8119: color = 12'h000;
            8120: color = 12'h000;
            8121: color = 12'h000;
            8122: color = 12'h000;
            8123: color = 12'hFFF;
            8124: color = 12'hFFF;
            8125: color = 12'hFFF;
            8126: color = 12'h000;
            8127: color = 12'h000;
            8128: color = 12'h000;
            8129: color = 12'h000;
            8130: color = 12'h000;
            8131: color = 12'h000;
            8132: color = 12'h000;
            8133: color = 12'h000;
            8134: color = 12'h000;
            8135: color = 12'h000;
            8136: color = 12'h000;
            8137: color = 12'h000;
            8138: color = 12'h000;
            8139: color = 12'h888;
            8140: color = 12'hFFF;
            8141: color = 12'hFFF;
            8142: color = 12'h777;
            8143: color = 12'h000;
            8144: color = 12'h000;
            8145: color = 12'h000;
            8146: color = 12'h000;
            8147: color = 12'h000;
            8148: color = 12'h000;
            8149: color = 12'h000;
            8150: color = 12'hFFF;
            8151: color = 12'hFFF;
            8152: color = 12'hFFF;
            8153: color = 12'h000;
            8154: color = 12'h000;
            8155: color = 12'h000;
            8156: color = 12'hFFF;
            8157: color = 12'hFFF;
            8158: color = 12'hFFF;
            8159: color = 12'h000;
            8160: color = 12'h000;
            8161: color = 12'h000;
            8162: color = 12'h000;
            8163: color = 12'h888;
            8164: color = 12'hFFF;
            8165: color = 12'hFFF;
            8166: color = 12'hFFF;
            8167: color = 12'hFFF;
            8168: color = 12'hFFF;
            8169: color = 12'hFFF;
            8170: color = 12'hFFF;
            8171: color = 12'hFFF;
            8172: color = 12'hCCC;
            8173: color = 12'h888;
            8174: color = 12'h888;
            8175: color = 12'h444;
            8176: color = 12'h000;
            8177: color = 12'hFFF;
            8178: color = 12'hFFF;
            8179: color = 12'hFFF;
            8180: color = 12'h000;
            8181: color = 12'h000;
            8182: color = 12'h000;
            8183: color = 12'h000;
            8184: color = 12'h000;
            8185: color = 12'h000;
            8186: color = 12'h000;
            8187: color = 12'h000;
            8188: color = 12'h000;
            8189: color = 12'h000;
            8190: color = 12'h000;
            8191: color = 12'h000;
            8192: color = 12'h000;
            8193: color = 12'h000;
            8194: color = 12'h000;
            8195: color = 12'h000;
            8196: color = 12'h000;
            8197: color = 12'h000;
            8198: color = 12'hFFF;
            8199: color = 12'hFFF;
            8200: color = 12'hFFF;
            8201: color = 12'h000;
            8202: color = 12'h000;
            8203: color = 12'h000;
            8204: color = 12'h000;
            8205: color = 12'h888;
            8206: color = 12'hFFF;
            8207: color = 12'hFFF;
            8208: color = 12'h777;
            8209: color = 12'h000;
            8210: color = 12'h000;
            8211: color = 12'h000;
            8212: color = 12'h000;
            8213: color = 12'h000;
            8214: color = 12'h888;
            8215: color = 12'hFFF;
            8216: color = 12'hFFF;
            8217: color = 12'h777;
            8218: color = 12'h000;
            8219: color = 12'h000;
            8220: color = 12'h000;
            8221: color = 12'h000;
            8222: color = 12'h000;
            8223: color = 12'h000;
            8224: color = 12'h000;
            8225: color = 12'h000;
            8226: color = 12'h000;
            8227: color = 12'h000;
            8228: color = 12'h000;
            8229: color = 12'h000;
            8230: color = 12'h000;
            8231: color = 12'h000;
            8232: color = 12'h000;
            8233: color = 12'h000;
            8234: color = 12'h000;
            8235: color = 12'h000;
            8236: color = 12'h000;
            8237: color = 12'hFFF;
            8238: color = 12'hFFF;
            8239: color = 12'hFFF;
            8240: color = 12'h000;
            8241: color = 12'h000;
            8242: color = 12'h000;
            8243: color = 12'hFFF;
            8244: color = 12'hFFF;
            8245: color = 12'hFFF;
            8246: color = 12'h000;
            8247: color = 12'h000;
            8248: color = 12'h000;
            8249: color = 12'h000;
            8250: color = 12'h000;
            8251: color = 12'h000;
            8252: color = 12'h000;
            8253: color = 12'h888;
            8254: color = 12'hFFF;
            8255: color = 12'hFFF;
            8256: color = 12'hFFF;
            8257: color = 12'hFFF;
            8258: color = 12'hFFF;
            8259: color = 12'hFFF;
            8260: color = 12'hFFF;
            8261: color = 12'hFFF;
            8262: color = 12'hFFF;
            8263: color = 12'hFFF;
            8264: color = 12'h000;
            8265: color = 12'h888;
            8266: color = 12'hFFF;
            8267: color = 12'hFFF;
            8268: color = 12'h777;
            8269: color = 12'h000;
            8270: color = 12'h000;
            8271: color = 12'h000;
            8272: color = 12'h000;
            8273: color = 12'h000;
            8274: color = 12'h000;
            8275: color = 12'h000;
            8276: color = 12'h000;
            8277: color = 12'h000;
            8278: color = 12'h000;
            8279: color = 12'hFFF;
            8280: color = 12'hFFF;
            8281: color = 12'hFFF;
            8282: color = 12'h000;
            8283: color = 12'h000;
            8284: color = 12'h000;
            8285: color = 12'h000;
            8286: color = 12'h000;
            8287: color = 12'h000;
            8288: color = 12'h000;
            8289: color = 12'h000;
            8290: color = 12'h000;
            8291: color = 12'h000;
            8292: color = 12'h000;
            8293: color = 12'h000;
            8294: color = 12'h000;
            8295: color = 12'h000;
            8296: color = 12'h000;
            8297: color = 12'h000;
            8298: color = 12'h000;
            8299: color = 12'h000;
            8300: color = 12'h000;
            8301: color = 12'h000;
            8302: color = 12'h000;
            8303: color = 12'h000;
            8304: color = 12'h000;
            8305: color = 12'h000;
            8306: color = 12'h000;
            8307: color = 12'h000;
            8308: color = 12'h000;
            8309: color = 12'h000;
            8310: color = 12'h000;
            8311: color = 12'h000;
            8312: color = 12'h000;
            8313: color = 12'h000;
            8314: color = 12'h000;
            8315: color = 12'h000;
            8316: color = 12'h000;
            8317: color = 12'h000;
            8318: color = 12'h000;
            8319: color = 12'h000;
            8320: color = 12'h000;
            8321: color = 12'h000;
            8322: color = 12'h000;
            8323: color = 12'h000;
            8324: color = 12'h000;
            8325: color = 12'h000;
            8326: color = 12'h000;
            8327: color = 12'h000;
            8328: color = 12'h000;
            8329: color = 12'h000;
            8330: color = 12'h000;
            8331: color = 12'h000;
            8332: color = 12'h000;
            8333: color = 12'h000;
            8334: color = 12'h000;
            8335: color = 12'h000;
            8336: color = 12'h000;
            8337: color = 12'h000;
            8338: color = 12'h000;
            8339: color = 12'h000;
            8340: color = 12'h000;
            8341: color = 12'h000;
            8342: color = 12'h000;
            8343: color = 12'h000;
            8344: color = 12'h000;
            8345: color = 12'h000;
            8346: color = 12'h000;
            8347: color = 12'h000;
            8348: color = 12'h000;
            8349: color = 12'h000;
            8350: color = 12'h000;
            8351: color = 12'h000;
            8352: color = 12'h000;
            8353: color = 12'h000;
            8354: color = 12'h000;
            8355: color = 12'h000;
            8356: color = 12'h000;
            8357: color = 12'h000;
            8358: color = 12'h000;
            8359: color = 12'h000;
            8360: color = 12'h000;
            8361: color = 12'h000;
            8362: color = 12'h000;
            8363: color = 12'h000;
            8364: color = 12'h000;
            8365: color = 12'h000;
            8366: color = 12'h000;
            8367: color = 12'h000;
            8368: color = 12'h000;
            8369: color = 12'h888;
            8370: color = 12'hFFF;
            8371: color = 12'hFFF;
            8372: color = 12'h777;
            8373: color = 12'h000;
            8374: color = 12'h000;
            8375: color = 12'h000;
            8376: color = 12'h000;
            8377: color = 12'h000;
            8378: color = 12'h000;
            8379: color = 12'h000;
            8380: color = 12'h000;
            8381: color = 12'h000;
            8382: color = 12'h000;
            8383: color = 12'h000;
            8384: color = 12'h000;
            8385: color = 12'h000;
            8386: color = 12'hFFF;
            8387: color = 12'hFFF;
            8388: color = 12'hFFF;
            8389: color = 12'h000;
            8390: color = 12'h000;
            8391: color = 12'h000;
            8392: color = 12'h000;
            8393: color = 12'h000;
            8394: color = 12'h000;
            8395: color = 12'h000;
            8396: color = 12'h000;
            8397: color = 12'h000;
            8398: color = 12'hFFF;
            8399: color = 12'hFFF;
            8400: color = 12'hFFF;
            8401: color = 12'hFFF;
            8402: color = 12'hFFF;
            8403: color = 12'hFFF;
            8404: color = 12'hFFF;
            8405: color = 12'hFFF;
            8406: color = 12'hEEE;
            8407: color = 12'h000;
            8408: color = 12'h000;
            8409: color = 12'h000;
            8410: color = 12'h000;
            8411: color = 12'h000;
            8412: color = 12'h000;
            8413: color = 12'h000;
            8414: color = 12'h777;
            8415: color = 12'hFFF;
            8416: color = 12'hFFF;
            8417: color = 12'hFFF;
            8418: color = 12'hEEE;
            8419: color = 12'h111;
            8420: color = 12'h000;
            8421: color = 12'h000;
            8422: color = 12'h000;
            8423: color = 12'h000;
            8424: color = 12'h000;
            8425: color = 12'h000;
            8426: color = 12'h777;
            8427: color = 12'hFFF;
            8428: color = 12'hFFF;
            8429: color = 12'hFFF;
            8430: color = 12'hEEE;
            8431: color = 12'h111;
            8432: color = 12'h000;
            8433: color = 12'h000;
            8434: color = 12'h000;
            8435: color = 12'h000;
            8436: color = 12'h000;
            8437: color = 12'h000;
            8438: color = 12'h000;
            8439: color = 12'h000;
            8440: color = 12'h000;
            8441: color = 12'h000;
            8442: color = 12'h000;
            8443: color = 12'hFFF;
            8444: color = 12'hFFF;
            8445: color = 12'hFFF;
            8446: color = 12'h000;
            8447: color = 12'h000;
            8448: color = 12'h000;
            8449: color = 12'h000;
            8450: color = 12'h000;
            8451: color = 12'h000;
            8452: color = 12'h000;
            8453: color = 12'h000;
            8454: color = 12'h000;
            8455: color = 12'h000;
            8456: color = 12'h000;
            8457: color = 12'h000;
            8458: color = 12'h000;
            8459: color = 12'h888;
            8460: color = 12'hFFF;
            8461: color = 12'hFFF;
            8462: color = 12'h777;
            8463: color = 12'h000;
            8464: color = 12'h000;
            8465: color = 12'h000;
            8466: color = 12'h000;
            8467: color = 12'h000;
            8468: color = 12'h000;
            8469: color = 12'h000;
            8470: color = 12'hFFF;
            8471: color = 12'hFFF;
            8472: color = 12'hFFF;
            8473: color = 12'h000;
            8474: color = 12'h000;
            8475: color = 12'h000;
            8476: color = 12'hFFF;
            8477: color = 12'hFFF;
            8478: color = 12'hFFF;
            8479: color = 12'h000;
            8480: color = 12'h000;
            8481: color = 12'h000;
            8482: color = 12'h000;
            8483: color = 12'h888;
            8484: color = 12'hFFF;
            8485: color = 12'hFFF;
            8486: color = 12'hFFF;
            8487: color = 12'hFFF;
            8488: color = 12'hFFF;
            8489: color = 12'hFFF;
            8490: color = 12'hFFF;
            8491: color = 12'hFFF;
            8492: color = 12'h777;
            8493: color = 12'h000;
            8494: color = 12'h000;
            8495: color = 12'h000;
            8496: color = 12'h000;
            8497: color = 12'hFFF;
            8498: color = 12'hFFF;
            8499: color = 12'hFFF;
            8500: color = 12'h000;
            8501: color = 12'h000;
            8502: color = 12'h000;
            8503: color = 12'h000;
            8504: color = 12'h000;
            8505: color = 12'h000;
            8506: color = 12'h000;
            8507: color = 12'h000;
            8508: color = 12'h000;
            8509: color = 12'h000;
            8510: color = 12'h000;
            8511: color = 12'h000;
            8512: color = 12'h000;
            8513: color = 12'h000;
            8514: color = 12'h000;
            8515: color = 12'h000;
            8516: color = 12'h000;
            8517: color = 12'h000;
            8518: color = 12'hFFF;
            8519: color = 12'hFFF;
            8520: color = 12'hFFF;
            8521: color = 12'h000;
            8522: color = 12'h000;
            8523: color = 12'h000;
            8524: color = 12'h000;
            8525: color = 12'h888;
            8526: color = 12'hFFF;
            8527: color = 12'hFFF;
            8528: color = 12'h777;
            8529: color = 12'h000;
            8530: color = 12'h000;
            8531: color = 12'h000;
            8532: color = 12'h000;
            8533: color = 12'h000;
            8534: color = 12'h888;
            8535: color = 12'hFFF;
            8536: color = 12'hFFF;
            8537: color = 12'h777;
            8538: color = 12'h000;
            8539: color = 12'h000;
            8540: color = 12'h000;
            8541: color = 12'h000;
            8542: color = 12'h000;
            8543: color = 12'h000;
            8544: color = 12'h000;
            8545: color = 12'h000;
            8546: color = 12'h000;
            8547: color = 12'h000;
            8548: color = 12'h000;
            8549: color = 12'h000;
            8550: color = 12'h000;
            8551: color = 12'h000;
            8552: color = 12'h000;
            8553: color = 12'h000;
            8554: color = 12'h000;
            8555: color = 12'h000;
            8556: color = 12'h000;
            8557: color = 12'hFFF;
            8558: color = 12'hFFF;
            8559: color = 12'hFFF;
            8560: color = 12'h000;
            8561: color = 12'h000;
            8562: color = 12'h000;
            8563: color = 12'hFFF;
            8564: color = 12'hFFF;
            8565: color = 12'hFFF;
            8566: color = 12'h000;
            8567: color = 12'h000;
            8568: color = 12'h000;
            8569: color = 12'h000;
            8570: color = 12'h000;
            8571: color = 12'h000;
            8572: color = 12'h000;
            8573: color = 12'h888;
            8574: color = 12'hFFF;
            8575: color = 12'hFFF;
            8576: color = 12'hFFF;
            8577: color = 12'hFFF;
            8578: color = 12'hFFF;
            8579: color = 12'hFFF;
            8580: color = 12'hFFF;
            8581: color = 12'hFFF;
            8582: color = 12'hFFF;
            8583: color = 12'hFFF;
            8584: color = 12'h000;
            8585: color = 12'h888;
            8586: color = 12'hFFF;
            8587: color = 12'hFFF;
            8588: color = 12'h777;
            8589: color = 12'h000;
            8590: color = 12'h000;
            8591: color = 12'h000;
            8592: color = 12'h000;
            8593: color = 12'h000;
            8594: color = 12'h000;
            8595: color = 12'h000;
            8596: color = 12'h000;
            8597: color = 12'h000;
            8598: color = 12'h000;
            8599: color = 12'hFFF;
            8600: color = 12'hFFF;
            8601: color = 12'hFFF;
            8602: color = 12'h000;
            8603: color = 12'h000;
            8604: color = 12'h000;
            8605: color = 12'h000;
            8606: color = 12'h000;
            8607: color = 12'h000;
            8608: color = 12'h000;
            8609: color = 12'h000;
            8610: color = 12'h000;
            8611: color = 12'h000;
            8612: color = 12'h000;
            8613: color = 12'h000;
            8614: color = 12'h000;
            8615: color = 12'h000;
            8616: color = 12'h000;
            8617: color = 12'h000;
            8618: color = 12'h000;
            8619: color = 12'h000;
            8620: color = 12'h000;
            8621: color = 12'h000;
            8622: color = 12'h000;
            8623: color = 12'h000;
            8624: color = 12'h000;
            8625: color = 12'h000;
            8626: color = 12'h000;
            8627: color = 12'h000;
            8628: color = 12'h000;
            8629: color = 12'h000;
            8630: color = 12'h000;
            8631: color = 12'h000;
            8632: color = 12'h000;
            8633: color = 12'h000;
            8634: color = 12'h000;
            8635: color = 12'h000;
            8636: color = 12'h000;
            8637: color = 12'h000;
            8638: color = 12'h000;
            8639: color = 12'h000;
            8640: color = 12'h000;
            8641: color = 12'h000;
            8642: color = 12'h000;
            8643: color = 12'h000;
            8644: color = 12'h000;
            8645: color = 12'h000;
            8646: color = 12'h000;
            8647: color = 12'h000;
            8648: color = 12'h000;
            8649: color = 12'h000;
            8650: color = 12'h000;
            8651: color = 12'h000;
            8652: color = 12'h000;
            8653: color = 12'h000;
            8654: color = 12'h000;
            8655: color = 12'h000;
            8656: color = 12'h000;
            8657: color = 12'h000;
            8658: color = 12'h000;
            8659: color = 12'h000;
            8660: color = 12'h000;
            8661: color = 12'h000;
            8662: color = 12'h000;
            8663: color = 12'h000;
            8664: color = 12'h000;
            8665: color = 12'h000;
            8666: color = 12'h000;
            8667: color = 12'h000;
            8668: color = 12'h000;
            8669: color = 12'h000;
            8670: color = 12'h000;
            8671: color = 12'h000;
            8672: color = 12'h000;
            8673: color = 12'h000;
            8674: color = 12'h000;
            8675: color = 12'h000;
            8676: color = 12'h000;
            8677: color = 12'h000;
            8678: color = 12'h000;
            8679: color = 12'h000;
            8680: color = 12'h000;
            8681: color = 12'h000;
            8682: color = 12'h000;
            8683: color = 12'h000;
            8684: color = 12'h000;
            8685: color = 12'h000;
            8686: color = 12'h000;
            8687: color = 12'h000;
            8688: color = 12'h000;
            8689: color = 12'h888;
            8690: color = 12'hFFF;
            8691: color = 12'hFFF;
            8692: color = 12'h777;
            8693: color = 12'h000;
            8694: color = 12'h000;
            8695: color = 12'h000;
            8696: color = 12'h000;
            8697: color = 12'h000;
            8698: color = 12'h000;
            8699: color = 12'h000;
            8700: color = 12'h000;
            8701: color = 12'h000;
            8702: color = 12'h000;
            8703: color = 12'h000;
            8704: color = 12'h000;
            8705: color = 12'h000;
            8706: color = 12'hFFF;
            8707: color = 12'hFFF;
            8708: color = 12'hFFF;
            8709: color = 12'h000;
            8710: color = 12'h000;
            8711: color = 12'h000;
            8712: color = 12'h000;
            8713: color = 12'h000;
            8714: color = 12'h000;
            8715: color = 12'h000;
            8716: color = 12'h000;
            8717: color = 12'h000;
            8718: color = 12'hFFF;
            8719: color = 12'hFFF;
            8720: color = 12'hFFF;
            8721: color = 12'h111;
            8722: color = 12'h000;
            8723: color = 12'h000;
            8724: color = 12'h000;
            8725: color = 12'h000;
            8726: color = 12'h000;
            8727: color = 12'h000;
            8728: color = 12'h000;
            8729: color = 12'h000;
            8730: color = 12'h000;
            8731: color = 12'h000;
            8732: color = 12'h000;
            8733: color = 12'h000;
            8734: color = 12'h000;
            8735: color = 12'h000;
            8736: color = 12'h000;
            8737: color = 12'h000;
            8738: color = 12'h111;
            8739: color = 12'hEEE;
            8740: color = 12'hFFF;
            8741: color = 12'hEEE;
            8742: color = 12'h000;
            8743: color = 12'h000;
            8744: color = 12'h000;
            8745: color = 12'h000;
            8746: color = 12'h000;
            8747: color = 12'h000;
            8748: color = 12'h000;
            8749: color = 12'h000;
            8750: color = 12'h111;
            8751: color = 12'hEEE;
            8752: color = 12'hFFF;
            8753: color = 12'hEEE;
            8754: color = 12'h000;
            8755: color = 12'h000;
            8756: color = 12'h000;
            8757: color = 12'h000;
            8758: color = 12'h000;
            8759: color = 12'h000;
            8760: color = 12'h000;
            8761: color = 12'h000;
            8762: color = 12'h000;
            8763: color = 12'hFFF;
            8764: color = 12'hFFF;
            8765: color = 12'hFFF;
            8766: color = 12'h000;
            8767: color = 12'h000;
            8768: color = 12'h000;
            8769: color = 12'h000;
            8770: color = 12'h000;
            8771: color = 12'h000;
            8772: color = 12'h000;
            8773: color = 12'h000;
            8774: color = 12'h000;
            8775: color = 12'h000;
            8776: color = 12'h000;
            8777: color = 12'h000;
            8778: color = 12'h000;
            8779: color = 12'h888;
            8780: color = 12'hFFF;
            8781: color = 12'hFFF;
            8782: color = 12'h777;
            8783: color = 12'h000;
            8784: color = 12'h000;
            8785: color = 12'h000;
            8786: color = 12'h000;
            8787: color = 12'h000;
            8788: color = 12'h000;
            8789: color = 12'h000;
            8790: color = 12'hFFF;
            8791: color = 12'hFFF;
            8792: color = 12'hFFF;
            8793: color = 12'h000;
            8794: color = 12'h000;
            8795: color = 12'h000;
            8796: color = 12'hFFF;
            8797: color = 12'hFFF;
            8798: color = 12'hFFF;
            8799: color = 12'h000;
            8800: color = 12'h000;
            8801: color = 12'h000;
            8802: color = 12'h000;
            8803: color = 12'h888;
            8804: color = 12'hFFF;
            8805: color = 12'hFFF;
            8806: color = 12'h888;
            8807: color = 12'h000;
            8808: color = 12'h000;
            8809: color = 12'h000;
            8810: color = 12'h000;
            8811: color = 12'h000;
            8812: color = 12'h000;
            8813: color = 12'h000;
            8814: color = 12'h000;
            8815: color = 12'h000;
            8816: color = 12'h000;
            8817: color = 12'hFFF;
            8818: color = 12'hFFF;
            8819: color = 12'hFFF;
            8820: color = 12'h000;
            8821: color = 12'h000;
            8822: color = 12'h000;
            8823: color = 12'h000;
            8824: color = 12'h000;
            8825: color = 12'h000;
            8826: color = 12'h000;
            8827: color = 12'h000;
            8828: color = 12'h000;
            8829: color = 12'h000;
            8830: color = 12'h000;
            8831: color = 12'h000;
            8832: color = 12'h000;
            8833: color = 12'h000;
            8834: color = 12'h000;
            8835: color = 12'h000;
            8836: color = 12'h000;
            8837: color = 12'h000;
            8838: color = 12'hFFF;
            8839: color = 12'hFFF;
            8840: color = 12'hFFF;
            8841: color = 12'h000;
            8842: color = 12'h000;
            8843: color = 12'h000;
            8844: color = 12'h000;
            8845: color = 12'h888;
            8846: color = 12'hFFF;
            8847: color = 12'hFFF;
            8848: color = 12'h777;
            8849: color = 12'h000;
            8850: color = 12'h000;
            8851: color = 12'h000;
            8852: color = 12'h000;
            8853: color = 12'h000;
            8854: color = 12'h888;
            8855: color = 12'hFFF;
            8856: color = 12'hFFF;
            8857: color = 12'h777;
            8858: color = 12'h000;
            8859: color = 12'h000;
            8860: color = 12'h000;
            8861: color = 12'h000;
            8862: color = 12'h000;
            8863: color = 12'h000;
            8864: color = 12'h000;
            8865: color = 12'h000;
            8866: color = 12'h000;
            8867: color = 12'h000;
            8868: color = 12'h000;
            8869: color = 12'h000;
            8870: color = 12'h000;
            8871: color = 12'h000;
            8872: color = 12'h000;
            8873: color = 12'h000;
            8874: color = 12'h000;
            8875: color = 12'h000;
            8876: color = 12'h000;
            8877: color = 12'hFFF;
            8878: color = 12'hFFF;
            8879: color = 12'hFFF;
            8880: color = 12'h000;
            8881: color = 12'h000;
            8882: color = 12'h000;
            8883: color = 12'hFFF;
            8884: color = 12'hFFF;
            8885: color = 12'hFFF;
            8886: color = 12'h000;
            8887: color = 12'h000;
            8888: color = 12'h000;
            8889: color = 12'h000;
            8890: color = 12'h777;
            8891: color = 12'hFFF;
            8892: color = 12'hFFF;
            8893: color = 12'h888;
            8894: color = 12'h000;
            8895: color = 12'h000;
            8896: color = 12'h000;
            8897: color = 12'h000;
            8898: color = 12'h000;
            8899: color = 12'h000;
            8900: color = 12'h111;
            8901: color = 12'hFFF;
            8902: color = 12'hFFF;
            8903: color = 12'hFFF;
            8904: color = 12'h000;
            8905: color = 12'h888;
            8906: color = 12'hFFF;
            8907: color = 12'hFFF;
            8908: color = 12'h777;
            8909: color = 12'h000;
            8910: color = 12'h000;
            8911: color = 12'h000;
            8912: color = 12'h000;
            8913: color = 12'h000;
            8914: color = 12'h000;
            8915: color = 12'h000;
            8916: color = 12'h000;
            8917: color = 12'h000;
            8918: color = 12'h000;
            8919: color = 12'hFFF;
            8920: color = 12'hFFF;
            8921: color = 12'hFFF;
            8922: color = 12'h000;
            8923: color = 12'h000;
            8924: color = 12'h000;
            8925: color = 12'h000;
            8926: color = 12'h000;
            8927: color = 12'h000;
            8928: color = 12'h000;
            8929: color = 12'h000;
            8930: color = 12'h000;
            8931: color = 12'h000;
            8932: color = 12'h000;
            8933: color = 12'h000;
            8934: color = 12'h000;
            8935: color = 12'h000;
            8936: color = 12'h000;
            8937: color = 12'h000;
            8938: color = 12'h000;
            8939: color = 12'h000;
            8940: color = 12'h000;
            8941: color = 12'h000;
            8942: color = 12'h000;
            8943: color = 12'h000;
            8944: color = 12'h000;
            8945: color = 12'h000;
            8946: color = 12'h000;
            8947: color = 12'h000;
            8948: color = 12'h000;
            8949: color = 12'h000;
            8950: color = 12'h000;
            8951: color = 12'h000;
            8952: color = 12'h000;
            8953: color = 12'h000;
            8954: color = 12'h000;
            8955: color = 12'h000;
            8956: color = 12'h000;
            8957: color = 12'h000;
            8958: color = 12'h000;
            8959: color = 12'h000;
            8960: color = 12'h000;
            8961: color = 12'h000;
            8962: color = 12'h000;
            8963: color = 12'h000;
            8964: color = 12'h000;
            8965: color = 12'h000;
            8966: color = 12'h000;
            8967: color = 12'h000;
            8968: color = 12'h000;
            8969: color = 12'h000;
            8970: color = 12'h000;
            8971: color = 12'h000;
            8972: color = 12'h000;
            8973: color = 12'h000;
            8974: color = 12'h000;
            8975: color = 12'h000;
            8976: color = 12'h000;
            8977: color = 12'h000;
            8978: color = 12'h000;
            8979: color = 12'h000;
            8980: color = 12'h000;
            8981: color = 12'h000;
            8982: color = 12'h000;
            8983: color = 12'h000;
            8984: color = 12'h000;
            8985: color = 12'h000;
            8986: color = 12'h000;
            8987: color = 12'h000;
            8988: color = 12'h000;
            8989: color = 12'h000;
            8990: color = 12'h000;
            8991: color = 12'h000;
            8992: color = 12'h000;
            8993: color = 12'h000;
            8994: color = 12'h000;
            8995: color = 12'h000;
            8996: color = 12'h000;
            8997: color = 12'h000;
            8998: color = 12'h000;
            8999: color = 12'h000;
            9000: color = 12'h000;
            9001: color = 12'h000;
            9002: color = 12'h000;
            9003: color = 12'h000;
            9004: color = 12'h000;
            9005: color = 12'h000;
            9006: color = 12'h000;
            9007: color = 12'h000;
            9008: color = 12'h000;
            9009: color = 12'h888;
            9010: color = 12'hFFF;
            9011: color = 12'hFFF;
            9012: color = 12'h777;
            9013: color = 12'h000;
            9014: color = 12'h000;
            9015: color = 12'h000;
            9016: color = 12'h000;
            9017: color = 12'h000;
            9018: color = 12'h000;
            9019: color = 12'h000;
            9020: color = 12'h000;
            9021: color = 12'h000;
            9022: color = 12'h000;
            9023: color = 12'h000;
            9024: color = 12'h000;
            9025: color = 12'h000;
            9026: color = 12'hFFF;
            9027: color = 12'hFFF;
            9028: color = 12'hFFF;
            9029: color = 12'h000;
            9030: color = 12'h000;
            9031: color = 12'h000;
            9032: color = 12'h000;
            9033: color = 12'h000;
            9034: color = 12'h000;
            9035: color = 12'h000;
            9036: color = 12'h000;
            9037: color = 12'h000;
            9038: color = 12'hFFF;
            9039: color = 12'hFFF;
            9040: color = 12'hFFF;
            9041: color = 12'h000;
            9042: color = 12'h000;
            9043: color = 12'h000;
            9044: color = 12'h000;
            9045: color = 12'h000;
            9046: color = 12'h000;
            9047: color = 12'h777;
            9048: color = 12'h888;
            9049: color = 12'h777;
            9050: color = 12'h000;
            9051: color = 12'h000;
            9052: color = 12'h000;
            9053: color = 12'h000;
            9054: color = 12'h000;
            9055: color = 12'h000;
            9056: color = 12'h000;
            9057: color = 12'h000;
            9058: color = 12'h000;
            9059: color = 12'hFFF;
            9060: color = 12'hFFF;
            9061: color = 12'hFFF;
            9062: color = 12'h000;
            9063: color = 12'h000;
            9064: color = 12'h000;
            9065: color = 12'h000;
            9066: color = 12'h000;
            9067: color = 12'h000;
            9068: color = 12'h000;
            9069: color = 12'h000;
            9070: color = 12'h000;
            9071: color = 12'hFFF;
            9072: color = 12'hFFF;
            9073: color = 12'hFFF;
            9074: color = 12'h000;
            9075: color = 12'h000;
            9076: color = 12'h000;
            9077: color = 12'h000;
            9078: color = 12'h000;
            9079: color = 12'h000;
            9080: color = 12'h000;
            9081: color = 12'h000;
            9082: color = 12'h000;
            9083: color = 12'hFFF;
            9084: color = 12'hFFF;
            9085: color = 12'hFFF;
            9086: color = 12'h000;
            9087: color = 12'h000;
            9088: color = 12'h000;
            9089: color = 12'h000;
            9090: color = 12'h000;
            9091: color = 12'h000;
            9092: color = 12'h000;
            9093: color = 12'h000;
            9094: color = 12'h000;
            9095: color = 12'h000;
            9096: color = 12'h000;
            9097: color = 12'h000;
            9098: color = 12'h000;
            9099: color = 12'h888;
            9100: color = 12'hFFF;
            9101: color = 12'hFFF;
            9102: color = 12'h777;
            9103: color = 12'h000;
            9104: color = 12'h000;
            9105: color = 12'h000;
            9106: color = 12'h000;
            9107: color = 12'h000;
            9108: color = 12'h000;
            9109: color = 12'h000;
            9110: color = 12'hFFF;
            9111: color = 12'hFFF;
            9112: color = 12'hFFF;
            9113: color = 12'h000;
            9114: color = 12'h000;
            9115: color = 12'h000;
            9116: color = 12'hFFF;
            9117: color = 12'hFFF;
            9118: color = 12'hFFF;
            9119: color = 12'h000;
            9120: color = 12'h000;
            9121: color = 12'h000;
            9122: color = 12'h000;
            9123: color = 12'h888;
            9124: color = 12'hFFF;
            9125: color = 12'hFFF;
            9126: color = 12'h777;
            9127: color = 12'h000;
            9128: color = 12'h000;
            9129: color = 12'h000;
            9130: color = 12'h000;
            9131: color = 12'h000;
            9132: color = 12'h444;
            9133: color = 12'h888;
            9134: color = 12'h888;
            9135: color = 12'h444;
            9136: color = 12'h000;
            9137: color = 12'hFFF;
            9138: color = 12'hFFF;
            9139: color = 12'hFFF;
            9140: color = 12'h000;
            9141: color = 12'h000;
            9142: color = 12'h000;
            9143: color = 12'h000;
            9144: color = 12'h000;
            9145: color = 12'h000;
            9146: color = 12'h000;
            9147: color = 12'h000;
            9148: color = 12'h000;
            9149: color = 12'h000;
            9150: color = 12'h000;
            9151: color = 12'h000;
            9152: color = 12'h000;
            9153: color = 12'h000;
            9154: color = 12'h000;
            9155: color = 12'h000;
            9156: color = 12'h000;
            9157: color = 12'h000;
            9158: color = 12'hFFF;
            9159: color = 12'hFFF;
            9160: color = 12'hFFF;
            9161: color = 12'h000;
            9162: color = 12'h000;
            9163: color = 12'h000;
            9164: color = 12'h000;
            9165: color = 12'h888;
            9166: color = 12'hFFF;
            9167: color = 12'hFFF;
            9168: color = 12'h777;
            9169: color = 12'h000;
            9170: color = 12'h000;
            9171: color = 12'h000;
            9172: color = 12'h000;
            9173: color = 12'h000;
            9174: color = 12'h888;
            9175: color = 12'hFFF;
            9176: color = 12'hFFF;
            9177: color = 12'h777;
            9178: color = 12'h000;
            9179: color = 12'h000;
            9180: color = 12'h000;
            9181: color = 12'h000;
            9182: color = 12'h000;
            9183: color = 12'h000;
            9184: color = 12'h000;
            9185: color = 12'h000;
            9186: color = 12'h000;
            9187: color = 12'h000;
            9188: color = 12'h000;
            9189: color = 12'h000;
            9190: color = 12'h000;
            9191: color = 12'h000;
            9192: color = 12'h000;
            9193: color = 12'h000;
            9194: color = 12'h000;
            9195: color = 12'h000;
            9196: color = 12'h000;
            9197: color = 12'hFFF;
            9198: color = 12'hFFF;
            9199: color = 12'hFFF;
            9200: color = 12'h000;
            9201: color = 12'h000;
            9202: color = 12'h000;
            9203: color = 12'hFFF;
            9204: color = 12'hFFF;
            9205: color = 12'hFFF;
            9206: color = 12'h000;
            9207: color = 12'h000;
            9208: color = 12'h000;
            9209: color = 12'h000;
            9210: color = 12'h888;
            9211: color = 12'hFFF;
            9212: color = 12'hFFF;
            9213: color = 12'h777;
            9214: color = 12'h000;
            9215: color = 12'h000;
            9216: color = 12'h000;
            9217: color = 12'h000;
            9218: color = 12'h000;
            9219: color = 12'h000;
            9220: color = 12'h000;
            9221: color = 12'hFFF;
            9222: color = 12'hFFF;
            9223: color = 12'hFFF;
            9224: color = 12'h000;
            9225: color = 12'h888;
            9226: color = 12'hFFF;
            9227: color = 12'hFFF;
            9228: color = 12'h777;
            9229: color = 12'h000;
            9230: color = 12'h000;
            9231: color = 12'h000;
            9232: color = 12'h000;
            9233: color = 12'h000;
            9234: color = 12'h000;
            9235: color = 12'h000;
            9236: color = 12'h000;
            9237: color = 12'h000;
            9238: color = 12'h000;
            9239: color = 12'hFFF;
            9240: color = 12'hFFF;
            9241: color = 12'hFFF;
            9242: color = 12'h000;
            9243: color = 12'h000;
            9244: color = 12'h000;
            9245: color = 12'h000;
            9246: color = 12'h000;
            9247: color = 12'h000;
            9248: color = 12'h000;
            9249: color = 12'h000;
            9250: color = 12'h000;
            9251: color = 12'h000;
            9252: color = 12'h000;
            9253: color = 12'h000;
            9254: color = 12'h000;
            9255: color = 12'h000;
            9256: color = 12'h000;
            9257: color = 12'h000;
            9258: color = 12'h000;
            9259: color = 12'h000;
            9260: color = 12'h000;
            9261: color = 12'h000;
            9262: color = 12'h000;
            9263: color = 12'h000;
            9264: color = 12'h000;
            9265: color = 12'h000;
            9266: color = 12'h000;
            9267: color = 12'h000;
            9268: color = 12'h000;
            9269: color = 12'h000;
            9270: color = 12'h000;
            9271: color = 12'h000;
            9272: color = 12'h000;
            9273: color = 12'h000;
            9274: color = 12'h000;
            9275: color = 12'h000;
            9276: color = 12'h000;
            9277: color = 12'h000;
            9278: color = 12'h000;
            9279: color = 12'h000;
            9280: color = 12'h000;
            9281: color = 12'h000;
            9282: color = 12'h000;
            9283: color = 12'h000;
            9284: color = 12'h000;
            9285: color = 12'h000;
            9286: color = 12'h000;
            9287: color = 12'h000;
            9288: color = 12'h000;
            9289: color = 12'h000;
            9290: color = 12'h000;
            9291: color = 12'h000;
            9292: color = 12'h000;
            9293: color = 12'h000;
            9294: color = 12'h000;
            9295: color = 12'h000;
            9296: color = 12'h000;
            9297: color = 12'h000;
            9298: color = 12'h000;
            9299: color = 12'h000;
            9300: color = 12'h000;
            9301: color = 12'h000;
            9302: color = 12'h000;
            9303: color = 12'h000;
            9304: color = 12'h000;
            9305: color = 12'h000;
            9306: color = 12'h000;
            9307: color = 12'h000;
            9308: color = 12'h000;
            9309: color = 12'h000;
            9310: color = 12'h000;
            9311: color = 12'h000;
            9312: color = 12'h000;
            9313: color = 12'h000;
            9314: color = 12'h000;
            9315: color = 12'h000;
            9316: color = 12'h000;
            9317: color = 12'h000;
            9318: color = 12'h000;
            9319: color = 12'h000;
            9320: color = 12'h000;
            9321: color = 12'h000;
            9322: color = 12'h000;
            9323: color = 12'h000;
            9324: color = 12'h000;
            9325: color = 12'h000;
            9326: color = 12'h000;
            9327: color = 12'h000;
            9328: color = 12'h000;
            9329: color = 12'h888;
            9330: color = 12'hFFF;
            9331: color = 12'hFFF;
            9332: color = 12'h777;
            9333: color = 12'h000;
            9334: color = 12'h000;
            9335: color = 12'h000;
            9336: color = 12'h000;
            9337: color = 12'h000;
            9338: color = 12'h000;
            9339: color = 12'h000;
            9340: color = 12'h000;
            9341: color = 12'h000;
            9342: color = 12'h000;
            9343: color = 12'h000;
            9344: color = 12'h000;
            9345: color = 12'h000;
            9346: color = 12'hFFF;
            9347: color = 12'hFFF;
            9348: color = 12'hFFF;
            9349: color = 12'h000;
            9350: color = 12'h000;
            9351: color = 12'h000;
            9352: color = 12'h000;
            9353: color = 12'h000;
            9354: color = 12'h000;
            9355: color = 12'h000;
            9356: color = 12'h000;
            9357: color = 12'h000;
            9358: color = 12'hEEE;
            9359: color = 12'hFFF;
            9360: color = 12'hEEE;
            9361: color = 12'h111;
            9362: color = 12'h000;
            9363: color = 12'h000;
            9364: color = 12'h000;
            9365: color = 12'h000;
            9366: color = 12'h111;
            9367: color = 12'hFFF;
            9368: color = 12'hFFF;
            9369: color = 12'hFFF;
            9370: color = 12'h000;
            9371: color = 12'h000;
            9372: color = 12'h000;
            9373: color = 12'h000;
            9374: color = 12'h000;
            9375: color = 12'h000;
            9376: color = 12'h000;
            9377: color = 12'h000;
            9378: color = 12'h111;
            9379: color = 12'hEEE;
            9380: color = 12'hFFF;
            9381: color = 12'hEEE;
            9382: color = 12'h000;
            9383: color = 12'h000;
            9384: color = 12'h000;
            9385: color = 12'h000;
            9386: color = 12'h000;
            9387: color = 12'h000;
            9388: color = 12'h000;
            9389: color = 12'h000;
            9390: color = 12'h111;
            9391: color = 12'hEEE;
            9392: color = 12'hFFF;
            9393: color = 12'hEEE;
            9394: color = 12'h000;
            9395: color = 12'h000;
            9396: color = 12'h000;
            9397: color = 12'h000;
            9398: color = 12'h000;
            9399: color = 12'h000;
            9400: color = 12'h000;
            9401: color = 12'h000;
            9402: color = 12'h000;
            9403: color = 12'hFFF;
            9404: color = 12'hFFF;
            9405: color = 12'hFFF;
            9406: color = 12'h111;
            9407: color = 12'h000;
            9408: color = 12'h000;
            9409: color = 12'h000;
            9410: color = 12'h000;
            9411: color = 12'h000;
            9412: color = 12'h000;
            9413: color = 12'h000;
            9414: color = 12'h000;
            9415: color = 12'h000;
            9416: color = 12'h000;
            9417: color = 12'h000;
            9418: color = 12'h000;
            9419: color = 12'h888;
            9420: color = 12'hFFF;
            9421: color = 12'hFFF;
            9422: color = 12'h777;
            9423: color = 12'h000;
            9424: color = 12'h000;
            9425: color = 12'h000;
            9426: color = 12'h000;
            9427: color = 12'h000;
            9428: color = 12'h000;
            9429: color = 12'h000;
            9430: color = 12'hFFF;
            9431: color = 12'hFFF;
            9432: color = 12'hFFF;
            9433: color = 12'h000;
            9434: color = 12'h000;
            9435: color = 12'h000;
            9436: color = 12'hEEE;
            9437: color = 12'hFFF;
            9438: color = 12'hEEE;
            9439: color = 12'h111;
            9440: color = 12'h000;
            9441: color = 12'h000;
            9442: color = 12'h000;
            9443: color = 12'h777;
            9444: color = 12'hFFF;
            9445: color = 12'hFFF;
            9446: color = 12'h888;
            9447: color = 12'h000;
            9448: color = 12'h000;
            9449: color = 12'h000;
            9450: color = 12'h000;
            9451: color = 12'h000;
            9452: color = 12'h888;
            9453: color = 12'hFFF;
            9454: color = 12'hFFF;
            9455: color = 12'h777;
            9456: color = 12'h000;
            9457: color = 12'hFFF;
            9458: color = 12'hFFF;
            9459: color = 12'hFFF;
            9460: color = 12'h000;
            9461: color = 12'h000;
            9462: color = 12'h000;
            9463: color = 12'h000;
            9464: color = 12'h000;
            9465: color = 12'h000;
            9466: color = 12'h000;
            9467: color = 12'h000;
            9468: color = 12'h000;
            9469: color = 12'h000;
            9470: color = 12'h000;
            9471: color = 12'h000;
            9472: color = 12'h000;
            9473: color = 12'h000;
            9474: color = 12'h000;
            9475: color = 12'h000;
            9476: color = 12'h000;
            9477: color = 12'h000;
            9478: color = 12'hEEE;
            9479: color = 12'hFFF;
            9480: color = 12'hEEE;
            9481: color = 12'h111;
            9482: color = 12'h000;
            9483: color = 12'h000;
            9484: color = 12'h000;
            9485: color = 12'h777;
            9486: color = 12'hFFF;
            9487: color = 12'hFFF;
            9488: color = 12'h888;
            9489: color = 12'h000;
            9490: color = 12'h000;
            9491: color = 12'h000;
            9492: color = 12'h000;
            9493: color = 12'h000;
            9494: color = 12'h888;
            9495: color = 12'hFFF;
            9496: color = 12'hFFF;
            9497: color = 12'h777;
            9498: color = 12'h000;
            9499: color = 12'h000;
            9500: color = 12'h000;
            9501: color = 12'h000;
            9502: color = 12'h000;
            9503: color = 12'h000;
            9504: color = 12'h000;
            9505: color = 12'h000;
            9506: color = 12'h000;
            9507: color = 12'h000;
            9508: color = 12'h000;
            9509: color = 12'h000;
            9510: color = 12'h000;
            9511: color = 12'h000;
            9512: color = 12'h000;
            9513: color = 12'h000;
            9514: color = 12'h000;
            9515: color = 12'h000;
            9516: color = 12'h111;
            9517: color = 12'hEEE;
            9518: color = 12'hFFF;
            9519: color = 12'hEEE;
            9520: color = 12'h000;
            9521: color = 12'h000;
            9522: color = 12'h000;
            9523: color = 12'hEEE;
            9524: color = 12'hFFF;
            9525: color = 12'hEEE;
            9526: color = 12'h111;
            9527: color = 12'h000;
            9528: color = 12'h000;
            9529: color = 12'h000;
            9530: color = 12'h777;
            9531: color = 12'hFFF;
            9532: color = 12'hFFF;
            9533: color = 12'h888;
            9534: color = 12'h000;
            9535: color = 12'h000;
            9536: color = 12'h000;
            9537: color = 12'h000;
            9538: color = 12'h000;
            9539: color = 12'h000;
            9540: color = 12'h111;
            9541: color = 12'hFFF;
            9542: color = 12'hFFF;
            9543: color = 12'hFFF;
            9544: color = 12'h000;
            9545: color = 12'h888;
            9546: color = 12'hFFF;
            9547: color = 12'hFFF;
            9548: color = 12'h777;
            9549: color = 12'h000;
            9550: color = 12'h000;
            9551: color = 12'h000;
            9552: color = 12'h000;
            9553: color = 12'h000;
            9554: color = 12'h000;
            9555: color = 12'h000;
            9556: color = 12'h000;
            9557: color = 12'h000;
            9558: color = 12'h000;
            9559: color = 12'hEEE;
            9560: color = 12'hFFF;
            9561: color = 12'hEEE;
            9562: color = 12'h111;
            9563: color = 12'h000;
            9564: color = 12'h000;
            9565: color = 12'h000;
            9566: color = 12'h000;
            9567: color = 12'h000;
            9568: color = 12'h000;
            9569: color = 12'h000;
            9570: color = 12'h000;
            9571: color = 12'h000;
            9572: color = 12'h000;
            9573: color = 12'h000;
            9574: color = 12'h000;
            9575: color = 12'h000;
            9576: color = 12'h000;
            9577: color = 12'h000;
            9578: color = 12'h000;
            9579: color = 12'h000;
            9580: color = 12'h000;
            9581: color = 12'h000;
            9582: color = 12'h000;
            9583: color = 12'h000;
            9584: color = 12'h000;
            9585: color = 12'h000;
            9586: color = 12'h000;
            9587: color = 12'h000;
            9588: color = 12'h000;
            9589: color = 12'h000;
            9590: color = 12'h000;
            9591: color = 12'h000;
            9592: color = 12'h000;
            9593: color = 12'h000;
            9594: color = 12'h000;
            9595: color = 12'h000;
            9596: color = 12'h000;
            9597: color = 12'h000;
            9598: color = 12'h000;
            9599: color = 12'h000;
            9600: color = 12'h000;
            9601: color = 12'h000;
            9602: color = 12'h000;
            9603: color = 12'h000;
            9604: color = 12'h000;
            9605: color = 12'h000;
            9606: color = 12'h000;
            9607: color = 12'h000;
            9608: color = 12'h000;
            9609: color = 12'h000;
            9610: color = 12'h000;
            9611: color = 12'h000;
            9612: color = 12'h000;
            9613: color = 12'h000;
            9614: color = 12'h000;
            9615: color = 12'h000;
            9616: color = 12'h000;
            9617: color = 12'h000;
            9618: color = 12'h000;
            9619: color = 12'h000;
            9620: color = 12'h000;
            9621: color = 12'h000;
            9622: color = 12'h000;
            9623: color = 12'h000;
            9624: color = 12'h000;
            9625: color = 12'h000;
            9626: color = 12'h000;
            9627: color = 12'h000;
            9628: color = 12'h000;
            9629: color = 12'h000;
            9630: color = 12'h000;
            9631: color = 12'h000;
            9632: color = 12'h000;
            9633: color = 12'h000;
            9634: color = 12'h000;
            9635: color = 12'h000;
            9636: color = 12'h000;
            9637: color = 12'h000;
            9638: color = 12'h000;
            9639: color = 12'h000;
            9640: color = 12'h000;
            9641: color = 12'h000;
            9642: color = 12'h000;
            9643: color = 12'h000;
            9644: color = 12'h000;
            9645: color = 12'h000;
            9646: color = 12'h000;
            9647: color = 12'h000;
            9648: color = 12'h000;
            9649: color = 12'h888;
            9650: color = 12'hFFF;
            9651: color = 12'hFFF;
            9652: color = 12'h777;
            9653: color = 12'h000;
            9654: color = 12'h000;
            9655: color = 12'h000;
            9656: color = 12'h000;
            9657: color = 12'h000;
            9658: color = 12'h000;
            9659: color = 12'h000;
            9660: color = 12'h000;
            9661: color = 12'h000;
            9662: color = 12'h000;
            9663: color = 12'h000;
            9664: color = 12'h000;
            9665: color = 12'h000;
            9666: color = 12'hFFF;
            9667: color = 12'hFFF;
            9668: color = 12'hFFF;
            9669: color = 12'h000;
            9670: color = 12'h000;
            9671: color = 12'h000;
            9672: color = 12'h000;
            9673: color = 12'h000;
            9674: color = 12'h000;
            9675: color = 12'h000;
            9676: color = 12'h000;
            9677: color = 12'h000;
            9678: color = 12'h000;
            9679: color = 12'h000;
            9680: color = 12'h111;
            9681: color = 12'hEEE;
            9682: color = 12'hFFF;
            9683: color = 12'hFFF;
            9684: color = 12'hFFF;
            9685: color = 12'hFFF;
            9686: color = 12'hFFF;
            9687: color = 12'hFFF;
            9688: color = 12'hFFF;
            9689: color = 12'hFFF;
            9690: color = 12'h000;
            9691: color = 12'h777;
            9692: color = 12'hFFF;
            9693: color = 12'hFFF;
            9694: color = 12'hFFF;
            9695: color = 12'hFFF;
            9696: color = 12'hFFF;
            9697: color = 12'hFFF;
            9698: color = 12'hEEE;
            9699: color = 12'h111;
            9700: color = 12'h000;
            9701: color = 12'h000;
            9702: color = 12'h000;
            9703: color = 12'h777;
            9704: color = 12'hFFF;
            9705: color = 12'hFFF;
            9706: color = 12'hFFF;
            9707: color = 12'hFFF;
            9708: color = 12'hFFF;
            9709: color = 12'hFFF;
            9710: color = 12'hEEE;
            9711: color = 12'h111;
            9712: color = 12'h000;
            9713: color = 12'h000;
            9714: color = 12'h000;
            9715: color = 12'h000;
            9716: color = 12'h000;
            9717: color = 12'h000;
            9718: color = 12'h000;
            9719: color = 12'h000;
            9720: color = 12'h000;
            9721: color = 12'h000;
            9722: color = 12'h000;
            9723: color = 12'hFFF;
            9724: color = 12'hFFF;
            9725: color = 12'hFFF;
            9726: color = 12'hFFF;
            9727: color = 12'hFFF;
            9728: color = 12'hFFF;
            9729: color = 12'hFFF;
            9730: color = 12'hFFF;
            9731: color = 12'hFFF;
            9732: color = 12'hFFF;
            9733: color = 12'hFFF;
            9734: color = 12'hFFF;
            9735: color = 12'hFFF;
            9736: color = 12'hFFF;
            9737: color = 12'hEEE;
            9738: color = 12'h000;
            9739: color = 12'h888;
            9740: color = 12'hFFF;
            9741: color = 12'hFFF;
            9742: color = 12'h777;
            9743: color = 12'h000;
            9744: color = 12'h000;
            9745: color = 12'h000;
            9746: color = 12'h000;
            9747: color = 12'h000;
            9748: color = 12'h000;
            9749: color = 12'h000;
            9750: color = 12'hFFF;
            9751: color = 12'hFFF;
            9752: color = 12'hFFF;
            9753: color = 12'h000;
            9754: color = 12'h000;
            9755: color = 12'h000;
            9756: color = 12'h000;
            9757: color = 12'h000;
            9758: color = 12'h111;
            9759: color = 12'hEEE;
            9760: color = 12'hFFF;
            9761: color = 12'hEEE;
            9762: color = 12'h000;
            9763: color = 12'h000;
            9764: color = 12'h000;
            9765: color = 12'h000;
            9766: color = 12'h888;
            9767: color = 12'hFFF;
            9768: color = 12'hFFF;
            9769: color = 12'hFFF;
            9770: color = 12'hFFF;
            9771: color = 12'hFFF;
            9772: color = 12'hFFF;
            9773: color = 12'hFFF;
            9774: color = 12'hFFF;
            9775: color = 12'h777;
            9776: color = 12'h000;
            9777: color = 12'hFFF;
            9778: color = 12'hFFF;
            9779: color = 12'hFFF;
            9780: color = 12'h000;
            9781: color = 12'h000;
            9782: color = 12'h000;
            9783: color = 12'h000;
            9784: color = 12'h000;
            9785: color = 12'h000;
            9786: color = 12'h000;
            9787: color = 12'h000;
            9788: color = 12'h000;
            9789: color = 12'h000;
            9790: color = 12'h000;
            9791: color = 12'h000;
            9792: color = 12'h000;
            9793: color = 12'h000;
            9794: color = 12'h000;
            9795: color = 12'h000;
            9796: color = 12'h000;
            9797: color = 12'h000;
            9798: color = 12'h000;
            9799: color = 12'h000;
            9800: color = 12'h111;
            9801: color = 12'hEEE;
            9802: color = 12'hFFF;
            9803: color = 12'hEEE;
            9804: color = 12'h000;
            9805: color = 12'h000;
            9806: color = 12'h000;
            9807: color = 12'h000;
            9808: color = 12'h888;
            9809: color = 12'hFFF;
            9810: color = 12'hFFF;
            9811: color = 12'hFFF;
            9812: color = 12'hFFF;
            9813: color = 12'hFFF;
            9814: color = 12'h888;
            9815: color = 12'h000;
            9816: color = 12'h000;
            9817: color = 12'h000;
            9818: color = 12'h000;
            9819: color = 12'h000;
            9820: color = 12'h000;
            9821: color = 12'h000;
            9822: color = 12'h000;
            9823: color = 12'h000;
            9824: color = 12'h000;
            9825: color = 12'h000;
            9826: color = 12'h777;
            9827: color = 12'hFFF;
            9828: color = 12'hFFF;
            9829: color = 12'hFFF;
            9830: color = 12'hFFF;
            9831: color = 12'hFFF;
            9832: color = 12'hFFF;
            9833: color = 12'hFFF;
            9834: color = 12'hFFF;
            9835: color = 12'hFFF;
            9836: color = 12'hEEE;
            9837: color = 12'h111;
            9838: color = 12'h000;
            9839: color = 12'h000;
            9840: color = 12'h000;
            9841: color = 12'h000;
            9842: color = 12'h000;
            9843: color = 12'h000;
            9844: color = 12'h000;
            9845: color = 12'h111;
            9846: color = 12'hEEE;
            9847: color = 12'hFFF;
            9848: color = 12'hEEE;
            9849: color = 12'h000;
            9850: color = 12'h000;
            9851: color = 12'h000;
            9852: color = 12'h000;
            9853: color = 12'h888;
            9854: color = 12'hFFF;
            9855: color = 12'hFFF;
            9856: color = 12'hFFF;
            9857: color = 12'hFFF;
            9858: color = 12'hFFF;
            9859: color = 12'hFFF;
            9860: color = 12'hFFF;
            9861: color = 12'hFFF;
            9862: color = 12'hFFF;
            9863: color = 12'hFFF;
            9864: color = 12'h000;
            9865: color = 12'h888;
            9866: color = 12'hFFF;
            9867: color = 12'hFFF;
            9868: color = 12'h777;
            9869: color = 12'h000;
            9870: color = 12'h000;
            9871: color = 12'h000;
            9872: color = 12'h000;
            9873: color = 12'h000;
            9874: color = 12'h000;
            9875: color = 12'h000;
            9876: color = 12'h000;
            9877: color = 12'h000;
            9878: color = 12'h000;
            9879: color = 12'h000;
            9880: color = 12'h000;
            9881: color = 12'h111;
            9882: color = 12'hEEE;
            9883: color = 12'hFFF;
            9884: color = 12'hEEE;
            9885: color = 12'h000;
            9886: color = 12'h000;
            9887: color = 12'h000;
            9888: color = 12'h000;
            9889: color = 12'h000;
            9890: color = 12'h000;
            9891: color = 12'h000;
            9892: color = 12'h000;
            9893: color = 12'h000;
            9894: color = 12'h000;
            9895: color = 12'h000;
            9896: color = 12'h000;
            9897: color = 12'h000;
            9898: color = 12'h000;
            9899: color = 12'h000;
            9900: color = 12'h000;
            9901: color = 12'h000;
            9902: color = 12'h000;
            9903: color = 12'h000;
            9904: color = 12'h000;
            9905: color = 12'h000;
            9906: color = 12'h000;
            9907: color = 12'h000;
            9908: color = 12'h000;
            9909: color = 12'h000;
            9910: color = 12'h000;
            9911: color = 12'h000;
            9912: color = 12'h000;
            9913: color = 12'h000;
            9914: color = 12'h000;
            9915: color = 12'h000;
            9916: color = 12'h000;
            9917: color = 12'h000;
            9918: color = 12'h000;
            9919: color = 12'h000;
            9920: color = 12'h000;
            9921: color = 12'h000;
            9922: color = 12'h000;
            9923: color = 12'h000;
            9924: color = 12'h000;
            9925: color = 12'h000;
            9926: color = 12'h000;
            9927: color = 12'h000;
            9928: color = 12'h000;
            9929: color = 12'h000;
            9930: color = 12'h000;
            9931: color = 12'h000;
            9932: color = 12'h000;
            9933: color = 12'h000;
            9934: color = 12'h000;
            9935: color = 12'h000;
            9936: color = 12'h000;
            9937: color = 12'h000;
            9938: color = 12'h000;
            9939: color = 12'h000;
            9940: color = 12'h000;
            9941: color = 12'h000;
            9942: color = 12'h000;
            9943: color = 12'h000;
            9944: color = 12'h000;
            9945: color = 12'h000;
            9946: color = 12'h000;
            9947: color = 12'h000;
            9948: color = 12'h000;
            9949: color = 12'h000;
            9950: color = 12'h000;
            9951: color = 12'h000;
            9952: color = 12'h000;
            9953: color = 12'h000;
            9954: color = 12'h000;
            9955: color = 12'h000;
            9956: color = 12'h000;
            9957: color = 12'h000;
            9958: color = 12'h000;
            9959: color = 12'h000;
            9960: color = 12'h000;
            9961: color = 12'h000;
            9962: color = 12'h000;
            9963: color = 12'h000;
            9964: color = 12'h000;
            9965: color = 12'h000;
            9966: color = 12'h000;
            9967: color = 12'h000;
            9968: color = 12'h000;
            9969: color = 12'h888;
            9970: color = 12'hFFF;
            9971: color = 12'hFFF;
            9972: color = 12'h777;
            9973: color = 12'h000;
            9974: color = 12'h000;
            9975: color = 12'h000;
            9976: color = 12'h000;
            9977: color = 12'h000;
            9978: color = 12'h000;
            9979: color = 12'h000;
            9980: color = 12'h000;
            9981: color = 12'h000;
            9982: color = 12'h000;
            9983: color = 12'h000;
            9984: color = 12'h000;
            9985: color = 12'h000;
            9986: color = 12'hFFF;
            9987: color = 12'hFFF;
            9988: color = 12'hFFF;
            9989: color = 12'h000;
            9990: color = 12'h000;
            9991: color = 12'h000;
            9992: color = 12'h000;
            9993: color = 12'h000;
            9994: color = 12'h000;
            9995: color = 12'h000;
            9996: color = 12'h000;
            9997: color = 12'h000;
            9998: color = 12'h000;
            9999: color = 12'h000;
            10000: color = 12'h000;
            10001: color = 12'hFFF;
            10002: color = 12'hFFF;
            10003: color = 12'hFFF;
            10004: color = 12'hFFF;
            10005: color = 12'hFFF;
            10006: color = 12'hFFF;
            10007: color = 12'hFFF;
            10008: color = 12'hFFF;
            10009: color = 12'hFFF;
            10010: color = 12'h000;
            10011: color = 12'h888;
            10012: color = 12'hFFF;
            10013: color = 12'hFFF;
            10014: color = 12'hFFF;
            10015: color = 12'hFFF;
            10016: color = 12'hFFF;
            10017: color = 12'hFFF;
            10018: color = 12'hFFF;
            10019: color = 12'h000;
            10020: color = 12'h000;
            10021: color = 12'h000;
            10022: color = 12'h000;
            10023: color = 12'h888;
            10024: color = 12'hFFF;
            10025: color = 12'hFFF;
            10026: color = 12'hFFF;
            10027: color = 12'hFFF;
            10028: color = 12'hFFF;
            10029: color = 12'hFFF;
            10030: color = 12'hFFF;
            10031: color = 12'h000;
            10032: color = 12'h000;
            10033: color = 12'h000;
            10034: color = 12'h000;
            10035: color = 12'h000;
            10036: color = 12'h000;
            10037: color = 12'h000;
            10038: color = 12'h000;
            10039: color = 12'h000;
            10040: color = 12'h000;
            10041: color = 12'h000;
            10042: color = 12'h000;
            10043: color = 12'hFFF;
            10044: color = 12'hFFF;
            10045: color = 12'hFFF;
            10046: color = 12'hFFF;
            10047: color = 12'hFFF;
            10048: color = 12'hFFF;
            10049: color = 12'hFFF;
            10050: color = 12'hFFF;
            10051: color = 12'hFFF;
            10052: color = 12'hFFF;
            10053: color = 12'hFFF;
            10054: color = 12'hFFF;
            10055: color = 12'hFFF;
            10056: color = 12'hFFF;
            10057: color = 12'hFFF;
            10058: color = 12'h000;
            10059: color = 12'h888;
            10060: color = 12'hFFF;
            10061: color = 12'hFFF;
            10062: color = 12'h777;
            10063: color = 12'h000;
            10064: color = 12'h000;
            10065: color = 12'h000;
            10066: color = 12'h000;
            10067: color = 12'h000;
            10068: color = 12'h000;
            10069: color = 12'h000;
            10070: color = 12'hFFF;
            10071: color = 12'hFFF;
            10072: color = 12'hFFF;
            10073: color = 12'h000;
            10074: color = 12'h000;
            10075: color = 12'h000;
            10076: color = 12'h000;
            10077: color = 12'h000;
            10078: color = 12'h000;
            10079: color = 12'hFFF;
            10080: color = 12'hFFF;
            10081: color = 12'hFFF;
            10082: color = 12'h000;
            10083: color = 12'h000;
            10084: color = 12'h000;
            10085: color = 12'h000;
            10086: color = 12'h888;
            10087: color = 12'hFFF;
            10088: color = 12'hFFF;
            10089: color = 12'hFFF;
            10090: color = 12'hFFF;
            10091: color = 12'hFFF;
            10092: color = 12'hFFF;
            10093: color = 12'hFFF;
            10094: color = 12'hFFF;
            10095: color = 12'h777;
            10096: color = 12'h000;
            10097: color = 12'hFFF;
            10098: color = 12'hFFF;
            10099: color = 12'hFFF;
            10100: color = 12'h000;
            10101: color = 12'h000;
            10102: color = 12'h000;
            10103: color = 12'h000;
            10104: color = 12'h000;
            10105: color = 12'h000;
            10106: color = 12'h000;
            10107: color = 12'h000;
            10108: color = 12'h000;
            10109: color = 12'h000;
            10110: color = 12'h000;
            10111: color = 12'h000;
            10112: color = 12'h000;
            10113: color = 12'h000;
            10114: color = 12'h000;
            10115: color = 12'h000;
            10116: color = 12'h000;
            10117: color = 12'h000;
            10118: color = 12'h000;
            10119: color = 12'h000;
            10120: color = 12'h000;
            10121: color = 12'hFFF;
            10122: color = 12'hFFF;
            10123: color = 12'hFFF;
            10124: color = 12'h000;
            10125: color = 12'h000;
            10126: color = 12'h000;
            10127: color = 12'h000;
            10128: color = 12'h888;
            10129: color = 12'hFFF;
            10130: color = 12'hFFF;
            10131: color = 12'hFFF;
            10132: color = 12'hFFF;
            10133: color = 12'hFFF;
            10134: color = 12'h777;
            10135: color = 12'h000;
            10136: color = 12'h000;
            10137: color = 12'h000;
            10138: color = 12'h000;
            10139: color = 12'h000;
            10140: color = 12'h000;
            10141: color = 12'h000;
            10142: color = 12'h000;
            10143: color = 12'h000;
            10144: color = 12'h000;
            10145: color = 12'h000;
            10146: color = 12'h888;
            10147: color = 12'hFFF;
            10148: color = 12'hFFF;
            10149: color = 12'hFFF;
            10150: color = 12'hFFF;
            10151: color = 12'hFFF;
            10152: color = 12'hFFF;
            10153: color = 12'hFFF;
            10154: color = 12'hFFF;
            10155: color = 12'hFFF;
            10156: color = 12'hFFF;
            10157: color = 12'h000;
            10158: color = 12'h000;
            10159: color = 12'h000;
            10160: color = 12'h000;
            10161: color = 12'h000;
            10162: color = 12'h000;
            10163: color = 12'h000;
            10164: color = 12'h000;
            10165: color = 12'h000;
            10166: color = 12'hFFF;
            10167: color = 12'hFFF;
            10168: color = 12'hFFF;
            10169: color = 12'h000;
            10170: color = 12'h000;
            10171: color = 12'h000;
            10172: color = 12'h000;
            10173: color = 12'h888;
            10174: color = 12'hFFF;
            10175: color = 12'hFFF;
            10176: color = 12'hFFF;
            10177: color = 12'hFFF;
            10178: color = 12'hFFF;
            10179: color = 12'hFFF;
            10180: color = 12'hFFF;
            10181: color = 12'hFFF;
            10182: color = 12'hFFF;
            10183: color = 12'hFFF;
            10184: color = 12'h000;
            10185: color = 12'h888;
            10186: color = 12'hFFF;
            10187: color = 12'hFFF;
            10188: color = 12'h777;
            10189: color = 12'h000;
            10190: color = 12'h000;
            10191: color = 12'h000;
            10192: color = 12'h000;
            10193: color = 12'h000;
            10194: color = 12'h000;
            10195: color = 12'h000;
            10196: color = 12'h000;
            10197: color = 12'h000;
            10198: color = 12'h000;
            10199: color = 12'h000;
            10200: color = 12'h000;
            10201: color = 12'h000;
            10202: color = 12'hFFF;
            10203: color = 12'hFFF;
            10204: color = 12'hFFF;
            10205: color = 12'h000;
            10206: color = 12'h000;
            10207: color = 12'h000;
            10208: color = 12'h000;
            10209: color = 12'h000;
            10210: color = 12'h000;
            10211: color = 12'h000;
            10212: color = 12'h000;
            10213: color = 12'h000;
            10214: color = 12'h000;
            10215: color = 12'h000;
            10216: color = 12'h000;
            10217: color = 12'h000;
            10218: color = 12'h000;
            10219: color = 12'h000;
            10220: color = 12'h000;
            10221: color = 12'h000;
            10222: color = 12'h000;
            10223: color = 12'h000;
            10224: color = 12'h000;
            10225: color = 12'h000;
            10226: color = 12'h000;
            10227: color = 12'h000;
            10228: color = 12'h000;
            10229: color = 12'h000;
            10230: color = 12'h000;
            10231: color = 12'h000;
            10232: color = 12'h000;
            10233: color = 12'h000;
            10234: color = 12'h000;
            10235: color = 12'h000;
            10236: color = 12'h000;
            10237: color = 12'h000;
            10238: color = 12'h000;
            10239: color = 12'h000;
            10240: color = 12'h000;
            10241: color = 12'h000;
            10242: color = 12'h000;
            10243: color = 12'h000;
            10244: color = 12'h000;
            10245: color = 12'h000;
            10246: color = 12'h000;
            10247: color = 12'h000;
            10248: color = 12'h000;
            10249: color = 12'h000;
            10250: color = 12'h000;
            10251: color = 12'h000;
            10252: color = 12'h000;
            10253: color = 12'h000;
            10254: color = 12'h000;
            10255: color = 12'h000;
            10256: color = 12'h000;
            10257: color = 12'h000;
            10258: color = 12'h000;
            10259: color = 12'h000;
            10260: color = 12'h000;
            10261: color = 12'h000;
            10262: color = 12'h000;
            10263: color = 12'h000;
            10264: color = 12'h000;
            10265: color = 12'h000;
            10266: color = 12'h000;
            10267: color = 12'h000;
            10268: color = 12'h000;
            10269: color = 12'h000;
            10270: color = 12'h000;
            10271: color = 12'h000;
            10272: color = 12'h000;
            10273: color = 12'h000;
            10274: color = 12'h000;
            10275: color = 12'h000;
            10276: color = 12'h000;
            10277: color = 12'h000;
            10278: color = 12'h000;
            10279: color = 12'h000;
            10280: color = 12'h000;
            10281: color = 12'h000;
            10282: color = 12'h000;
            10283: color = 12'h000;
            10284: color = 12'h000;
            10285: color = 12'h000;
            10286: color = 12'h000;
            10287: color = 12'h000;
            10288: color = 12'h000;
            10289: color = 12'h777;
            10290: color = 12'hFFF;
            10291: color = 12'hFFF;
            10292: color = 12'h777;
            10293: color = 12'h000;
            10294: color = 12'h000;
            10295: color = 12'h000;
            10296: color = 12'h000;
            10297: color = 12'h000;
            10298: color = 12'h000;
            10299: color = 12'h000;
            10300: color = 12'h000;
            10301: color = 12'h000;
            10302: color = 12'h000;
            10303: color = 12'h000;
            10304: color = 12'h000;
            10305: color = 12'h000;
            10306: color = 12'hEEE;
            10307: color = 12'hFFF;
            10308: color = 12'hEEE;
            10309: color = 12'h000;
            10310: color = 12'h000;
            10311: color = 12'h000;
            10312: color = 12'h000;
            10313: color = 12'h000;
            10314: color = 12'h000;
            10315: color = 12'h000;
            10316: color = 12'h000;
            10317: color = 12'h000;
            10318: color = 12'h000;
            10319: color = 12'h000;
            10320: color = 12'h000;
            10321: color = 12'hEEE;
            10322: color = 12'hFFF;
            10323: color = 12'hFFF;
            10324: color = 12'hFFF;
            10325: color = 12'hFFF;
            10326: color = 12'hFFF;
            10327: color = 12'hFFF;
            10328: color = 12'hFFF;
            10329: color = 12'hEEE;
            10330: color = 12'h000;
            10331: color = 12'h777;
            10332: color = 12'hFFF;
            10333: color = 12'hFFF;
            10334: color = 12'hFFF;
            10335: color = 12'hFFF;
            10336: color = 12'hFFF;
            10337: color = 12'hFFF;
            10338: color = 12'hEEE;
            10339: color = 12'h000;
            10340: color = 12'h000;
            10341: color = 12'h000;
            10342: color = 12'h000;
            10343: color = 12'h777;
            10344: color = 12'hFFF;
            10345: color = 12'hFFF;
            10346: color = 12'hFFF;
            10347: color = 12'hFFF;
            10348: color = 12'hFFF;
            10349: color = 12'hFFF;
            10350: color = 12'hEEE;
            10351: color = 12'h000;
            10352: color = 12'h000;
            10353: color = 12'h000;
            10354: color = 12'h000;
            10355: color = 12'h000;
            10356: color = 12'h000;
            10357: color = 12'h000;
            10358: color = 12'h000;
            10359: color = 12'h000;
            10360: color = 12'h000;
            10361: color = 12'h000;
            10362: color = 12'h000;
            10363: color = 12'hEEE;
            10364: color = 12'hFFF;
            10365: color = 12'hFFF;
            10366: color = 12'hFFF;
            10367: color = 12'hFFF;
            10368: color = 12'hFFF;
            10369: color = 12'hFFF;
            10370: color = 12'hFFF;
            10371: color = 12'hFFF;
            10372: color = 12'hFFF;
            10373: color = 12'hFFF;
            10374: color = 12'hFFF;
            10375: color = 12'hFFF;
            10376: color = 12'hFFF;
            10377: color = 12'hEEE;
            10378: color = 12'h000;
            10379: color = 12'h777;
            10380: color = 12'hFFF;
            10381: color = 12'hFFF;
            10382: color = 12'h777;
            10383: color = 12'h000;
            10384: color = 12'h000;
            10385: color = 12'h000;
            10386: color = 12'h000;
            10387: color = 12'h000;
            10388: color = 12'h000;
            10389: color = 12'h000;
            10390: color = 12'hEEE;
            10391: color = 12'hFFF;
            10392: color = 12'hEEE;
            10393: color = 12'h000;
            10394: color = 12'h000;
            10395: color = 12'h000;
            10396: color = 12'h000;
            10397: color = 12'h000;
            10398: color = 12'h000;
            10399: color = 12'hEEE;
            10400: color = 12'hFFF;
            10401: color = 12'hEEE;
            10402: color = 12'h000;
            10403: color = 12'h000;
            10404: color = 12'h000;
            10405: color = 12'h000;
            10406: color = 12'h777;
            10407: color = 12'hFFF;
            10408: color = 12'hFFF;
            10409: color = 12'hFFF;
            10410: color = 12'hFFF;
            10411: color = 12'hFFF;
            10412: color = 12'hFFF;
            10413: color = 12'hFFF;
            10414: color = 12'hFFF;
            10415: color = 12'h777;
            10416: color = 12'h000;
            10417: color = 12'hEEE;
            10418: color = 12'hFFF;
            10419: color = 12'hEEE;
            10420: color = 12'h000;
            10421: color = 12'h000;
            10422: color = 12'h000;
            10423: color = 12'h000;
            10424: color = 12'h000;
            10425: color = 12'h000;
            10426: color = 12'h000;
            10427: color = 12'h000;
            10428: color = 12'h000;
            10429: color = 12'h000;
            10430: color = 12'h000;
            10431: color = 12'h000;
            10432: color = 12'h000;
            10433: color = 12'h000;
            10434: color = 12'h000;
            10435: color = 12'h000;
            10436: color = 12'h000;
            10437: color = 12'h000;
            10438: color = 12'h000;
            10439: color = 12'h000;
            10440: color = 12'h000;
            10441: color = 12'hEEE;
            10442: color = 12'hFFF;
            10443: color = 12'hEEE;
            10444: color = 12'h000;
            10445: color = 12'h000;
            10446: color = 12'h000;
            10447: color = 12'h000;
            10448: color = 12'h777;
            10449: color = 12'hFFF;
            10450: color = 12'hFFF;
            10451: color = 12'hFFF;
            10452: color = 12'hFFF;
            10453: color = 12'hFFF;
            10454: color = 12'h777;
            10455: color = 12'h000;
            10456: color = 12'h000;
            10457: color = 12'h000;
            10458: color = 12'h000;
            10459: color = 12'h000;
            10460: color = 12'h000;
            10461: color = 12'h000;
            10462: color = 12'h000;
            10463: color = 12'h000;
            10464: color = 12'h000;
            10465: color = 12'h000;
            10466: color = 12'h777;
            10467: color = 12'hFFF;
            10468: color = 12'hFFF;
            10469: color = 12'hFFF;
            10470: color = 12'hFFF;
            10471: color = 12'hFFF;
            10472: color = 12'hFFF;
            10473: color = 12'hFFF;
            10474: color = 12'hFFF;
            10475: color = 12'hFFF;
            10476: color = 12'hEEE;
            10477: color = 12'h000;
            10478: color = 12'h000;
            10479: color = 12'h000;
            10480: color = 12'h000;
            10481: color = 12'h000;
            10482: color = 12'h000;
            10483: color = 12'h000;
            10484: color = 12'h000;
            10485: color = 12'h000;
            10486: color = 12'hEEE;
            10487: color = 12'hFFF;
            10488: color = 12'hEEE;
            10489: color = 12'h000;
            10490: color = 12'h000;
            10491: color = 12'h000;
            10492: color = 12'h000;
            10493: color = 12'h777;
            10494: color = 12'hFFF;
            10495: color = 12'hFFF;
            10496: color = 12'hFFF;
            10497: color = 12'hFFF;
            10498: color = 12'hFFF;
            10499: color = 12'hFFF;
            10500: color = 12'hFFF;
            10501: color = 12'hFFF;
            10502: color = 12'hFFF;
            10503: color = 12'hEEE;
            10504: color = 12'h000;
            10505: color = 12'h777;
            10506: color = 12'hFFF;
            10507: color = 12'hFFF;
            10508: color = 12'h777;
            10509: color = 12'h000;
            10510: color = 12'h000;
            10511: color = 12'h000;
            10512: color = 12'h000;
            10513: color = 12'h000;
            10514: color = 12'h000;
            10515: color = 12'h000;
            10516: color = 12'h000;
            10517: color = 12'h000;
            10518: color = 12'h000;
            10519: color = 12'h000;
            10520: color = 12'h000;
            10521: color = 12'h000;
            10522: color = 12'hEEE;
            10523: color = 12'hFFF;
            10524: color = 12'hEEE;
            10525: color = 12'h000;
            10526: color = 12'h000;
            10527: color = 12'h000;
            10528: color = 12'h000;
            10529: color = 12'h000;
            10530: color = 12'h000;
            10531: color = 12'h000;
            10532: color = 12'h000;
            10533: color = 12'h000;
            10534: color = 12'h000;
            10535: color = 12'h000;
            10536: color = 12'h000;
            10537: color = 12'h000;
            10538: color = 12'h000;
            10539: color = 12'h000;
            10540: color = 12'h000;
            10541: color = 12'h000;
            10542: color = 12'h000;
            10543: color = 12'h000;
            10544: color = 12'h000;
            10545: color = 12'h000;
            10546: color = 12'h000;
            10547: color = 12'h000;
            10548: color = 12'h000;
            10549: color = 12'h000;
            10550: color = 12'h000;
            10551: color = 12'h000;
            10552: color = 12'h000;
            10553: color = 12'h000;
            10554: color = 12'h000;
            10555: color = 12'h000;
            10556: color = 12'h000;
            10557: color = 12'h000;
            10558: color = 12'h000;
            10559: color = 12'h000;
            10560: color = 12'h000;
            10561: color = 12'h000;
            10562: color = 12'h000;
            10563: color = 12'h000;
            10564: color = 12'h000;
            10565: color = 12'h000;
            10566: color = 12'h000;
            10567: color = 12'h000;
            10568: color = 12'h000;
            10569: color = 12'h000;
            10570: color = 12'h000;
            10571: color = 12'h000;
            10572: color = 12'h000;
            10573: color = 12'h000;
            10574: color = 12'h000;
            10575: color = 12'h000;
            10576: color = 12'h000;
            10577: color = 12'h000;
            10578: color = 12'h000;
            10579: color = 12'h000;
            10580: color = 12'h000;
            10581: color = 12'h000;
            10582: color = 12'h000;
            10583: color = 12'h000;
            10584: color = 12'h000;
            10585: color = 12'h000;
            10586: color = 12'h000;
            10587: color = 12'h000;
            10588: color = 12'h000;
            10589: color = 12'h000;
            10590: color = 12'h000;
            10591: color = 12'h000;
            10592: color = 12'h000;
            10593: color = 12'h000;
            10594: color = 12'h000;
            10595: color = 12'h000;
            10596: color = 12'h000;
            10597: color = 12'h000;
            10598: color = 12'h000;
            10599: color = 12'h000;
            10600: color = 12'h000;
            10601: color = 12'h000;
            10602: color = 12'h000;
            10603: color = 12'h000;
            10604: color = 12'h000;
            10605: color = 12'h000;
            10606: color = 12'h000;
            10607: color = 12'h000;
            10608: color = 12'h000;
            10609: color = 12'h000;
            10610: color = 12'h000;
            10611: color = 12'h000;
            10612: color = 12'h000;
            10613: color = 12'h000;
            10614: color = 12'h000;
            10615: color = 12'h000;
            10616: color = 12'h000;
            10617: color = 12'h000;
            10618: color = 12'h000;
            10619: color = 12'h000;
            10620: color = 12'h000;
            10621: color = 12'h000;
            10622: color = 12'h000;
            10623: color = 12'h000;
            10624: color = 12'h000;
            10625: color = 12'h000;
            10626: color = 12'h000;
            10627: color = 12'h000;
            10628: color = 12'h000;
            10629: color = 12'h000;
            10630: color = 12'h000;
            10631: color = 12'h000;
            10632: color = 12'h000;
            10633: color = 12'h000;
            10634: color = 12'h000;
            10635: color = 12'h000;
            10636: color = 12'h000;
            10637: color = 12'h000;
            10638: color = 12'h000;
            10639: color = 12'h000;
            10640: color = 12'h000;
            10641: color = 12'h000;
            10642: color = 12'h000;
            10643: color = 12'h000;
            10644: color = 12'h000;
            10645: color = 12'h000;
            10646: color = 12'h000;
            10647: color = 12'h000;
            10648: color = 12'h000;
            10649: color = 12'h000;
            10650: color = 12'h000;
            10651: color = 12'h000;
            10652: color = 12'h000;
            10653: color = 12'h000;
            10654: color = 12'h000;
            10655: color = 12'h000;
            10656: color = 12'h000;
            10657: color = 12'h000;
            10658: color = 12'h000;
            10659: color = 12'h000;
            10660: color = 12'h000;
            10661: color = 12'h000;
            10662: color = 12'h000;
            10663: color = 12'h000;
            10664: color = 12'h000;
            10665: color = 12'h000;
            10666: color = 12'h000;
            10667: color = 12'h000;
            10668: color = 12'h000;
            10669: color = 12'h000;
            10670: color = 12'h000;
            10671: color = 12'h000;
            10672: color = 12'h000;
            10673: color = 12'h000;
            10674: color = 12'h000;
            10675: color = 12'h000;
            10676: color = 12'h000;
            10677: color = 12'h000;
            10678: color = 12'h000;
            10679: color = 12'h000;
            10680: color = 12'h000;
            10681: color = 12'h000;
            10682: color = 12'h000;
            10683: color = 12'h000;
            10684: color = 12'h000;
            10685: color = 12'h000;
            10686: color = 12'h000;
            10687: color = 12'h000;
            10688: color = 12'h000;
            10689: color = 12'h000;
            10690: color = 12'h000;
            10691: color = 12'h000;
            10692: color = 12'h000;
            10693: color = 12'h000;
            10694: color = 12'h000;
            10695: color = 12'h000;
            10696: color = 12'h000;
            10697: color = 12'h000;
            10698: color = 12'h000;
            10699: color = 12'h000;
            10700: color = 12'h000;
            10701: color = 12'h000;
            10702: color = 12'h000;
            10703: color = 12'h000;
            10704: color = 12'h000;
            10705: color = 12'h000;
            10706: color = 12'h000;
            10707: color = 12'h000;
            10708: color = 12'h000;
            10709: color = 12'h000;
            10710: color = 12'h000;
            10711: color = 12'h000;
            10712: color = 12'h000;
            10713: color = 12'h000;
            10714: color = 12'h000;
            10715: color = 12'h000;
            10716: color = 12'h000;
            10717: color = 12'h000;
            10718: color = 12'h000;
            10719: color = 12'h000;
            10720: color = 12'h000;
            10721: color = 12'h000;
            10722: color = 12'h000;
            10723: color = 12'h000;
            10724: color = 12'h000;
            10725: color = 12'h000;
            10726: color = 12'h000;
            10727: color = 12'h000;
            10728: color = 12'h000;
            10729: color = 12'h000;
            10730: color = 12'h000;
            10731: color = 12'h000;
            10732: color = 12'h000;
            10733: color = 12'h000;
            10734: color = 12'h000;
            10735: color = 12'h000;
            10736: color = 12'h000;
            10737: color = 12'h000;
            10738: color = 12'h000;
            10739: color = 12'h000;
            10740: color = 12'h000;
            10741: color = 12'h000;
            10742: color = 12'h000;
            10743: color = 12'h000;
            10744: color = 12'h000;
            10745: color = 12'h000;
            10746: color = 12'h000;
            10747: color = 12'h000;
            10748: color = 12'h000;
            10749: color = 12'h000;
            10750: color = 12'h000;
            10751: color = 12'h000;
            10752: color = 12'h000;
            10753: color = 12'h000;
            10754: color = 12'h000;
            10755: color = 12'h000;
            10756: color = 12'h000;
            10757: color = 12'h000;
            10758: color = 12'h000;
            10759: color = 12'h000;
            10760: color = 12'h000;
            10761: color = 12'h000;
            10762: color = 12'h000;
            10763: color = 12'h000;
            10764: color = 12'h000;
            10765: color = 12'h000;
            10766: color = 12'h000;
            10767: color = 12'h000;
            10768: color = 12'h000;
            10769: color = 12'h000;
            10770: color = 12'h000;
            10771: color = 12'h000;
            10772: color = 12'h000;
            10773: color = 12'h000;
            10774: color = 12'h000;
            10775: color = 12'h000;
            10776: color = 12'h000;
            10777: color = 12'h000;
            10778: color = 12'h000;
            10779: color = 12'h000;
            10780: color = 12'h000;
            10781: color = 12'h000;
            10782: color = 12'h000;
            10783: color = 12'h000;
            10784: color = 12'h000;
            10785: color = 12'h000;
            10786: color = 12'h000;
            10787: color = 12'h000;
            10788: color = 12'h000;
            10789: color = 12'h000;
            10790: color = 12'h000;
            10791: color = 12'h000;
            10792: color = 12'h000;
            10793: color = 12'h000;
            10794: color = 12'h000;
            10795: color = 12'h000;
            10796: color = 12'h000;
            10797: color = 12'h000;
            10798: color = 12'h000;
            10799: color = 12'h000;
            10800: color = 12'h000;
            10801: color = 12'h000;
            10802: color = 12'h000;
            10803: color = 12'h000;
            10804: color = 12'h000;
            10805: color = 12'h000;
            10806: color = 12'h000;
            10807: color = 12'h000;
            10808: color = 12'h000;
            10809: color = 12'h000;
            10810: color = 12'h000;
            10811: color = 12'h000;
            10812: color = 12'h000;
            10813: color = 12'h000;
            10814: color = 12'h000;
            10815: color = 12'h000;
            10816: color = 12'h000;
            10817: color = 12'h000;
            10818: color = 12'h000;
            10819: color = 12'h000;
            10820: color = 12'h000;
            10821: color = 12'h000;
            10822: color = 12'h000;
            10823: color = 12'h000;
            10824: color = 12'h000;
            10825: color = 12'h000;
            10826: color = 12'h000;
            10827: color = 12'h000;
            10828: color = 12'h000;
            10829: color = 12'h000;
            10830: color = 12'h000;
            10831: color = 12'h000;
            10832: color = 12'h000;
            10833: color = 12'h000;
            10834: color = 12'h000;
            10835: color = 12'h000;
            10836: color = 12'h000;
            10837: color = 12'h000;
            10838: color = 12'h000;
            10839: color = 12'h000;
            10840: color = 12'h000;
            10841: color = 12'h000;
            10842: color = 12'h000;
            10843: color = 12'h000;
            10844: color = 12'h000;
            10845: color = 12'h000;
            10846: color = 12'h000;
            10847: color = 12'h000;
            10848: color = 12'h000;
            10849: color = 12'h000;
            10850: color = 12'h000;
            10851: color = 12'h000;
            10852: color = 12'h000;
            10853: color = 12'h000;
            10854: color = 12'h000;
            10855: color = 12'h000;
            10856: color = 12'h000;
            10857: color = 12'h000;
            10858: color = 12'h000;
            10859: color = 12'h000;
            10860: color = 12'h000;
            10861: color = 12'h000;
            10862: color = 12'h000;
            10863: color = 12'h000;
            10864: color = 12'h000;
            10865: color = 12'h000;
            10866: color = 12'h000;
            10867: color = 12'h000;
            10868: color = 12'h000;
            10869: color = 12'h000;
            10870: color = 12'h000;
            10871: color = 12'h000;
            10872: color = 12'h000;
            10873: color = 12'h000;
            10874: color = 12'h000;
            10875: color = 12'h000;
            10876: color = 12'h000;
            10877: color = 12'h000;
            10878: color = 12'h000;
            10879: color = 12'h000;
            10880: color = 12'h000;
            10881: color = 12'h000;
            10882: color = 12'h000;
            10883: color = 12'h000;
            10884: color = 12'h000;
            10885: color = 12'h000;
            10886: color = 12'h000;
            10887: color = 12'h000;
            10888: color = 12'h000;
            10889: color = 12'h000;
            10890: color = 12'h000;
            10891: color = 12'h000;
            10892: color = 12'h000;
            10893: color = 12'h000;
            10894: color = 12'h000;
            10895: color = 12'h000;
            10896: color = 12'h000;
            10897: color = 12'h000;
            10898: color = 12'h000;
            10899: color = 12'h000;
            10900: color = 12'h000;
            10901: color = 12'h000;
            10902: color = 12'h000;
            10903: color = 12'h000;
            10904: color = 12'h000;
            10905: color = 12'h000;
            10906: color = 12'h000;
            10907: color = 12'h000;
            10908: color = 12'h000;
            10909: color = 12'h000;
            10910: color = 12'h000;
            10911: color = 12'h000;
            10912: color = 12'h000;
            10913: color = 12'h000;
            10914: color = 12'h000;
            10915: color = 12'h000;
            10916: color = 12'h000;
            10917: color = 12'h000;
            10918: color = 12'h000;
            10919: color = 12'h000;
            10920: color = 12'h000;
            10921: color = 12'h000;
            10922: color = 12'h000;
            10923: color = 12'h000;
            10924: color = 12'h000;
            10925: color = 12'h000;
            10926: color = 12'h000;
            10927: color = 12'h000;
            10928: color = 12'h000;
            10929: color = 12'h000;
            10930: color = 12'h000;
            10931: color = 12'h000;
            10932: color = 12'h000;
            10933: color = 12'h000;
            10934: color = 12'h000;
            10935: color = 12'h000;
            10936: color = 12'h000;
            10937: color = 12'h000;
            10938: color = 12'h000;
            10939: color = 12'h000;
            10940: color = 12'h000;
            10941: color = 12'h000;
            10942: color = 12'h000;
            10943: color = 12'h000;
            10944: color = 12'h000;
            10945: color = 12'h000;
            10946: color = 12'h000;
            10947: color = 12'h000;
            10948: color = 12'h000;
            10949: color = 12'h000;
            10950: color = 12'h000;
            10951: color = 12'h000;
            10952: color = 12'h000;
            10953: color = 12'h000;
            10954: color = 12'h000;
            10955: color = 12'h000;
            10956: color = 12'h000;
            10957: color = 12'h000;
            10958: color = 12'h000;
            10959: color = 12'h000;
            10960: color = 12'h000;
            10961: color = 12'h000;
            10962: color = 12'h000;
            10963: color = 12'h000;
            10964: color = 12'h000;
            10965: color = 12'h000;
            10966: color = 12'h000;
            10967: color = 12'h000;
            10968: color = 12'h000;
            10969: color = 12'h000;
            10970: color = 12'h000;
            10971: color = 12'h000;
            10972: color = 12'h000;
            10973: color = 12'h000;
            10974: color = 12'h000;
            10975: color = 12'h000;
            10976: color = 12'h000;
            10977: color = 12'h000;
            10978: color = 12'h000;
            10979: color = 12'h000;
            10980: color = 12'h000;
            10981: color = 12'h000;
            10982: color = 12'h000;
            10983: color = 12'h000;
            10984: color = 12'h000;
            10985: color = 12'h000;
            10986: color = 12'h000;
            10987: color = 12'h000;
            10988: color = 12'h000;
            10989: color = 12'h000;
            10990: color = 12'h000;
            10991: color = 12'h000;
            10992: color = 12'h000;
            10993: color = 12'h000;
            10994: color = 12'h000;
            10995: color = 12'h000;
            10996: color = 12'h000;
            10997: color = 12'h000;
            10998: color = 12'h000;
            10999: color = 12'h000;
            11000: color = 12'h000;
            11001: color = 12'h000;
            11002: color = 12'h000;
            11003: color = 12'h000;
            11004: color = 12'h000;
            11005: color = 12'h000;
            11006: color = 12'h000;
            11007: color = 12'h000;
            11008: color = 12'h000;
            11009: color = 12'h000;
            11010: color = 12'h000;
            11011: color = 12'h000;
            11012: color = 12'h000;
            11013: color = 12'h000;
            11014: color = 12'h000;
            11015: color = 12'h000;
            11016: color = 12'h000;
            11017: color = 12'h000;
            11018: color = 12'h000;
            11019: color = 12'h000;
            11020: color = 12'h000;
            11021: color = 12'h000;
            11022: color = 12'h000;
            11023: color = 12'h000;
            11024: color = 12'h000;
            11025: color = 12'h000;
            11026: color = 12'h000;
            11027: color = 12'h000;
            11028: color = 12'h000;
            11029: color = 12'h000;
            11030: color = 12'h000;
            11031: color = 12'h000;
            11032: color = 12'h000;
            11033: color = 12'h000;
            11034: color = 12'h000;
            11035: color = 12'h000;
            11036: color = 12'h000;
            11037: color = 12'h000;
            11038: color = 12'h000;
            11039: color = 12'h000;
            11040: color = 12'h000;
            11041: color = 12'h000;
            11042: color = 12'h000;
            11043: color = 12'h000;
            11044: color = 12'h000;
            11045: color = 12'h000;
            11046: color = 12'h000;
            11047: color = 12'h000;
            11048: color = 12'h000;
            11049: color = 12'h000;
            11050: color = 12'h000;
            11051: color = 12'h000;
            11052: color = 12'h000;
            11053: color = 12'h000;
            11054: color = 12'h000;
            11055: color = 12'h000;
            11056: color = 12'h000;
            11057: color = 12'h000;
            11058: color = 12'h000;
            11059: color = 12'h000;
            11060: color = 12'h000;
            11061: color = 12'h000;
            11062: color = 12'h000;
            11063: color = 12'h000;
            11064: color = 12'h000;
            11065: color = 12'h000;
            11066: color = 12'h000;
            11067: color = 12'h000;
            11068: color = 12'h000;
            11069: color = 12'h000;
            11070: color = 12'h000;
            11071: color = 12'h000;
            11072: color = 12'h000;
            11073: color = 12'h000;
            11074: color = 12'h000;
            11075: color = 12'h000;
            11076: color = 12'h000;
            11077: color = 12'h000;
            11078: color = 12'h000;
            11079: color = 12'h000;
            11080: color = 12'h000;
            11081: color = 12'h000;
            11082: color = 12'h000;
            11083: color = 12'h000;
            11084: color = 12'h000;
            11085: color = 12'h000;
            11086: color = 12'h000;
            11087: color = 12'h000;
            11088: color = 12'h000;
            11089: color = 12'h000;
            11090: color = 12'h000;
            11091: color = 12'h000;
            11092: color = 12'h000;
            11093: color = 12'h000;
            11094: color = 12'h000;
            11095: color = 12'h000;
            11096: color = 12'h000;
            11097: color = 12'h000;
            11098: color = 12'h000;
            11099: color = 12'h000;
            11100: color = 12'h000;
            11101: color = 12'h000;
            11102: color = 12'h000;
            11103: color = 12'h000;
            11104: color = 12'h000;
            11105: color = 12'h000;
            11106: color = 12'h000;
            11107: color = 12'h000;
            11108: color = 12'h000;
            11109: color = 12'h000;
            11110: color = 12'h000;
            11111: color = 12'h000;
            11112: color = 12'h000;
            11113: color = 12'h000;
            11114: color = 12'h000;
            11115: color = 12'h000;
            11116: color = 12'h000;
            11117: color = 12'h000;
            11118: color = 12'h000;
            11119: color = 12'h000;
            11120: color = 12'h000;
            11121: color = 12'h000;
            11122: color = 12'h000;
            11123: color = 12'h000;
            11124: color = 12'h000;
            11125: color = 12'h000;
            11126: color = 12'h000;
            11127: color = 12'h000;
            11128: color = 12'h000;
            11129: color = 12'h000;
            11130: color = 12'h000;
            11131: color = 12'h000;
            11132: color = 12'h000;
            11133: color = 12'h000;
            11134: color = 12'h000;
            11135: color = 12'h000;
            11136: color = 12'h000;
            11137: color = 12'h000;
            11138: color = 12'h000;
            11139: color = 12'h000;
            11140: color = 12'h000;
            11141: color = 12'h000;
            11142: color = 12'h000;
            11143: color = 12'h000;
            11144: color = 12'h000;
            11145: color = 12'h000;
            11146: color = 12'h000;
            11147: color = 12'h000;
            11148: color = 12'h000;
            11149: color = 12'h000;
            11150: color = 12'h000;
            11151: color = 12'h000;
            11152: color = 12'h000;
            11153: color = 12'h000;
            11154: color = 12'h000;
            11155: color = 12'h000;
            11156: color = 12'h000;
            11157: color = 12'h000;
            11158: color = 12'h000;
            11159: color = 12'h000;
            11160: color = 12'h000;
            11161: color = 12'h000;
            11162: color = 12'h000;
            11163: color = 12'h000;
            11164: color = 12'h000;
            11165: color = 12'h000;
            11166: color = 12'h000;
            11167: color = 12'h000;
            11168: color = 12'h000;
            11169: color = 12'h000;
            11170: color = 12'h000;
            11171: color = 12'h000;
            11172: color = 12'h000;
            11173: color = 12'h000;
            11174: color = 12'h000;
            11175: color = 12'h000;
            11176: color = 12'h000;
            11177: color = 12'h000;
            11178: color = 12'h000;
            11179: color = 12'h000;
            11180: color = 12'h000;
            11181: color = 12'h000;
            11182: color = 12'h000;
            11183: color = 12'h000;
            11184: color = 12'h000;
            11185: color = 12'h000;
            11186: color = 12'h000;
            11187: color = 12'h000;
            11188: color = 12'h000;
            11189: color = 12'h000;
            11190: color = 12'h000;
            11191: color = 12'h000;
            11192: color = 12'h000;
            11193: color = 12'h000;
            11194: color = 12'h000;
            11195: color = 12'h000;
            11196: color = 12'h000;
            11197: color = 12'h000;
            11198: color = 12'h000;
            11199: color = 12'h000;
            11200: color = 12'h000;
            11201: color = 12'h000;
            11202: color = 12'h000;
            11203: color = 12'h000;
            11204: color = 12'h000;
            11205: color = 12'h000;
            11206: color = 12'h000;
            11207: color = 12'h000;
            11208: color = 12'h000;
            11209: color = 12'h000;
            11210: color = 12'h000;
            11211: color = 12'h000;
            11212: color = 12'h000;
            11213: color = 12'h000;
            11214: color = 12'h000;
            11215: color = 12'h000;
            11216: color = 12'h000;
            11217: color = 12'h000;
            11218: color = 12'h000;
            11219: color = 12'h000;
            11220: color = 12'h000;
            11221: color = 12'h000;
            11222: color = 12'h000;
            11223: color = 12'h000;
            11224: color = 12'h000;
            11225: color = 12'h000;
            11226: color = 12'h000;
            11227: color = 12'h000;
            11228: color = 12'h000;
            11229: color = 12'h000;
            11230: color = 12'h000;
            11231: color = 12'h000;
            11232: color = 12'h000;
            11233: color = 12'h000;
            11234: color = 12'h000;
            11235: color = 12'h000;
            11236: color = 12'h000;
            11237: color = 12'h000;
            11238: color = 12'h000;
            11239: color = 12'h000;
            11240: color = 12'h000;
            11241: color = 12'h000;
            11242: color = 12'h000;
            11243: color = 12'h000;
            11244: color = 12'h000;
            11245: color = 12'h000;
            11246: color = 12'h000;
            11247: color = 12'h000;
            11248: color = 12'h000;
            11249: color = 12'h000;
            11250: color = 12'h000;
            11251: color = 12'h000;
            11252: color = 12'h000;
            11253: color = 12'h000;
            11254: color = 12'h000;
            11255: color = 12'h000;
            11256: color = 12'h000;
            11257: color = 12'h000;
            11258: color = 12'h000;
            11259: color = 12'h000;
            11260: color = 12'h000;
            11261: color = 12'h000;
            11262: color = 12'h000;
            11263: color = 12'h000;
            11264: color = 12'h000;
            11265: color = 12'h000;
            11266: color = 12'h000;
            11267: color = 12'h000;
            11268: color = 12'h000;
            11269: color = 12'h000;
            11270: color = 12'h000;
            11271: color = 12'h000;
            11272: color = 12'h000;
            11273: color = 12'h000;
            11274: color = 12'h000;
            11275: color = 12'h000;
            11276: color = 12'h000;
            11277: color = 12'h000;
            11278: color = 12'h000;
            11279: color = 12'h000;
            11280: color = 12'h000;
            11281: color = 12'h000;
            11282: color = 12'h000;
            11283: color = 12'h000;
            11284: color = 12'h000;
            11285: color = 12'h000;
            11286: color = 12'h000;
            11287: color = 12'h000;
            11288: color = 12'h000;
            11289: color = 12'h000;
            11290: color = 12'h000;
            11291: color = 12'h000;
            11292: color = 12'h000;
            11293: color = 12'h000;
            11294: color = 12'h000;
            11295: color = 12'h000;
            11296: color = 12'h000;
            11297: color = 12'h000;
            11298: color = 12'h000;
            11299: color = 12'h000;
            11300: color = 12'h000;
            11301: color = 12'h000;
            11302: color = 12'h000;
            11303: color = 12'h000;
            11304: color = 12'h000;
            11305: color = 12'h000;
            11306: color = 12'h000;
            11307: color = 12'h000;
            11308: color = 12'h000;
            11309: color = 12'h000;
            11310: color = 12'h000;
            11311: color = 12'h000;
            11312: color = 12'h000;
            11313: color = 12'h000;
            11314: color = 12'h000;
            11315: color = 12'h000;
            11316: color = 12'h000;
            11317: color = 12'h000;
            11318: color = 12'h000;
            11319: color = 12'h000;
            11320: color = 12'h000;
            11321: color = 12'h000;
            11322: color = 12'h000;
            11323: color = 12'h000;
            11324: color = 12'h000;
            11325: color = 12'h000;
            11326: color = 12'h000;
            11327: color = 12'h000;
            11328: color = 12'h000;
            11329: color = 12'h000;
            11330: color = 12'h000;
            11331: color = 12'h000;
            11332: color = 12'h000;
            11333: color = 12'h000;
            11334: color = 12'h000;
            11335: color = 12'h000;
            11336: color = 12'h000;
            11337: color = 12'h000;
            11338: color = 12'h000;
            11339: color = 12'h000;
            11340: color = 12'h000;
            11341: color = 12'h000;
            11342: color = 12'h000;
            11343: color = 12'h000;
            11344: color = 12'h000;
            11345: color = 12'h000;
            11346: color = 12'h000;
            11347: color = 12'h000;
            11348: color = 12'h000;
            11349: color = 12'h000;
            11350: color = 12'h000;
            11351: color = 12'h000;
            11352: color = 12'h000;
            11353: color = 12'h000;
            11354: color = 12'h000;
            11355: color = 12'h000;
            11356: color = 12'h000;
            11357: color = 12'h000;
            11358: color = 12'h000;
            11359: color = 12'h000;
            11360: color = 12'h000;
            11361: color = 12'h000;
            11362: color = 12'h000;
            11363: color = 12'h000;
            11364: color = 12'h000;
            11365: color = 12'h000;
            11366: color = 12'h000;
            11367: color = 12'h000;
            11368: color = 12'h000;
            11369: color = 12'h000;
            11370: color = 12'h000;
            11371: color = 12'h000;
            11372: color = 12'h000;
            11373: color = 12'h000;
            11374: color = 12'h000;
            11375: color = 12'h000;
            11376: color = 12'h000;
            11377: color = 12'h000;
            11378: color = 12'h000;
            11379: color = 12'h000;
            11380: color = 12'h000;
            11381: color = 12'h000;
            11382: color = 12'h000;
            11383: color = 12'h000;
            11384: color = 12'h000;
            11385: color = 12'h000;
            11386: color = 12'h000;
            11387: color = 12'h000;
            11388: color = 12'h000;
            11389: color = 12'h000;
            11390: color = 12'h000;
            11391: color = 12'h000;
            11392: color = 12'h000;
            11393: color = 12'h000;
            11394: color = 12'h000;
            11395: color = 12'h000;
            11396: color = 12'h000;
            11397: color = 12'h000;
            11398: color = 12'h000;
            11399: color = 12'h000;
            11400: color = 12'h000;
            11401: color = 12'h000;
            11402: color = 12'h000;
            11403: color = 12'h000;
            11404: color = 12'h000;
            11405: color = 12'h000;
            11406: color = 12'h000;
            11407: color = 12'h000;
            11408: color = 12'h000;
            11409: color = 12'h000;
            11410: color = 12'h000;
            11411: color = 12'h000;
            11412: color = 12'h000;
            11413: color = 12'h000;
            11414: color = 12'h000;
            11415: color = 12'h000;
            11416: color = 12'h000;
            11417: color = 12'h000;
            11418: color = 12'h000;
            11419: color = 12'h000;
            11420: color = 12'h000;
            11421: color = 12'h000;
            11422: color = 12'h000;
            11423: color = 12'h000;
            11424: color = 12'h000;
            11425: color = 12'h000;
            11426: color = 12'h000;
            11427: color = 12'h000;
            11428: color = 12'h000;
            11429: color = 12'h000;
            11430: color = 12'h000;
            11431: color = 12'h000;
            11432: color = 12'h000;
            11433: color = 12'h000;
            11434: color = 12'h000;
            11435: color = 12'h000;
            11436: color = 12'h000;
            11437: color = 12'h000;
            11438: color = 12'h000;
            11439: color = 12'h000;
            11440: color = 12'h000;
            11441: color = 12'h000;
            11442: color = 12'h000;
            11443: color = 12'h000;
            11444: color = 12'h000;
            11445: color = 12'h000;
            11446: color = 12'h000;
            11447: color = 12'h000;
            11448: color = 12'h000;
            11449: color = 12'h000;
            11450: color = 12'h000;
            11451: color = 12'h000;
            11452: color = 12'h000;
            11453: color = 12'h000;
            11454: color = 12'h000;
            11455: color = 12'h000;
            11456: color = 12'h000;
            11457: color = 12'h000;
            11458: color = 12'h000;
            11459: color = 12'h000;
            11460: color = 12'h000;
            11461: color = 12'h000;
            11462: color = 12'h000;
            11463: color = 12'h000;
            11464: color = 12'h000;
            11465: color = 12'h000;
            11466: color = 12'h000;
            11467: color = 12'h000;
            11468: color = 12'h000;
            11469: color = 12'h000;
            11470: color = 12'h000;
            11471: color = 12'h000;
            11472: color = 12'h000;
            11473: color = 12'h000;
            11474: color = 12'h000;
            11475: color = 12'h000;
            11476: color = 12'h000;
            11477: color = 12'h000;
            11478: color = 12'h000;
            11479: color = 12'h000;
            11480: color = 12'h000;
            11481: color = 12'h000;
            11482: color = 12'h000;
            11483: color = 12'h000;
            11484: color = 12'h000;
            11485: color = 12'h000;
            11486: color = 12'h000;
            11487: color = 12'h000;
            11488: color = 12'h000;
            11489: color = 12'h000;
            11490: color = 12'h000;
            11491: color = 12'h000;
            11492: color = 12'h000;
            11493: color = 12'h000;
            11494: color = 12'h000;
            11495: color = 12'h000;
            11496: color = 12'h000;
            11497: color = 12'h000;
            11498: color = 12'h000;
            11499: color = 12'h000;
            11500: color = 12'h000;
            11501: color = 12'h000;
            11502: color = 12'h000;
            11503: color = 12'h000;
            11504: color = 12'h000;
            11505: color = 12'h000;
            11506: color = 12'h000;
            11507: color = 12'h000;
            11508: color = 12'h000;
            11509: color = 12'h000;
            11510: color = 12'h000;
            11511: color = 12'h000;
            11512: color = 12'h000;
            11513: color = 12'h000;
            11514: color = 12'h000;
            11515: color = 12'h000;
            11516: color = 12'h000;
            11517: color = 12'h000;
            11518: color = 12'h000;
            11519: color = 12'h000;
            11520: color = 12'h000;
            11521: color = 12'h000;
            11522: color = 12'h000;
            11523: color = 12'h000;
            11524: color = 12'h000;
            11525: color = 12'h000;
            11526: color = 12'h000;
            11527: color = 12'h000;
            11528: color = 12'h000;
            11529: color = 12'h000;
            11530: color = 12'h000;
            11531: color = 12'h000;
            11532: color = 12'h000;
            11533: color = 12'h000;
            11534: color = 12'h000;
            11535: color = 12'h000;
            11536: color = 12'h000;
            11537: color = 12'h000;
            11538: color = 12'h000;
            11539: color = 12'h000;
            11540: color = 12'h000;
            11541: color = 12'h000;
            11542: color = 12'h000;
            11543: color = 12'h000;
            11544: color = 12'h000;
            11545: color = 12'h000;
            11546: color = 12'h000;
            11547: color = 12'h000;
            11548: color = 12'h000;
            11549: color = 12'h000;
            11550: color = 12'h000;
            11551: color = 12'h000;
            11552: color = 12'h000;
            11553: color = 12'h000;
            11554: color = 12'h000;
            11555: color = 12'h000;
            11556: color = 12'h000;
            11557: color = 12'h000;
            11558: color = 12'h000;
            11559: color = 12'h000;
            11560: color = 12'h000;
            11561: color = 12'h000;
            11562: color = 12'h000;
            11563: color = 12'h000;
            11564: color = 12'h000;
            11565: color = 12'h000;
            11566: color = 12'h000;
            11567: color = 12'h000;
            11568: color = 12'h000;
            11569: color = 12'h000;
            11570: color = 12'h000;
            11571: color = 12'h000;
            11572: color = 12'h000;
            11573: color = 12'h000;
            11574: color = 12'h000;
            11575: color = 12'h000;
            11576: color = 12'h000;
            11577: color = 12'h000;
            11578: color = 12'h000;
            11579: color = 12'h000;
            11580: color = 12'h000;
            11581: color = 12'h000;
            11582: color = 12'h000;
            11583: color = 12'h000;
            11584: color = 12'h000;
            11585: color = 12'h000;
            11586: color = 12'h000;
            11587: color = 12'h000;
            11588: color = 12'h000;
            11589: color = 12'h000;
            11590: color = 12'h000;
            11591: color = 12'h000;
            11592: color = 12'h000;
            11593: color = 12'h000;
            11594: color = 12'h000;
            11595: color = 12'h000;
            11596: color = 12'h000;
            11597: color = 12'h000;
            11598: color = 12'h000;
            11599: color = 12'h000;
            11600: color = 12'h000;
            11601: color = 12'h000;
            11602: color = 12'h000;
            11603: color = 12'h000;
            11604: color = 12'h000;
            11605: color = 12'h000;
            11606: color = 12'h000;
            11607: color = 12'h000;
            11608: color = 12'h000;
            11609: color = 12'h000;
            11610: color = 12'h000;
            11611: color = 12'h000;
            11612: color = 12'h000;
            11613: color = 12'h000;
            11614: color = 12'h000;
            11615: color = 12'h000;
            11616: color = 12'h000;
            11617: color = 12'h000;
            11618: color = 12'h000;
            11619: color = 12'h000;
            11620: color = 12'h000;
            11621: color = 12'h000;
            11622: color = 12'h000;
            11623: color = 12'h000;
            11624: color = 12'h000;
            11625: color = 12'h000;
            11626: color = 12'h000;
            11627: color = 12'h000;
            11628: color = 12'h000;
            11629: color = 12'h000;
            11630: color = 12'h000;
            11631: color = 12'h000;
            11632: color = 12'h000;
            11633: color = 12'h000;
            11634: color = 12'h000;
            11635: color = 12'h000;
            11636: color = 12'h000;
            11637: color = 12'h000;
            11638: color = 12'h000;
            11639: color = 12'h000;
            11640: color = 12'h000;
            11641: color = 12'h000;
            11642: color = 12'h000;
            11643: color = 12'h000;
            11644: color = 12'h000;
            11645: color = 12'h000;
            11646: color = 12'h000;
            11647: color = 12'h000;
            11648: color = 12'h000;
            11649: color = 12'h000;
            11650: color = 12'h000;
            11651: color = 12'h000;
            11652: color = 12'h000;
            11653: color = 12'h000;
            11654: color = 12'h000;
            11655: color = 12'h000;
            11656: color = 12'h000;
            11657: color = 12'h000;
            11658: color = 12'h000;
            11659: color = 12'h000;
            11660: color = 12'h000;
            11661: color = 12'h000;
            11662: color = 12'h000;
            11663: color = 12'h000;
            11664: color = 12'h000;
            11665: color = 12'h000;
            11666: color = 12'h000;
            11667: color = 12'h000;
            11668: color = 12'h000;
            11669: color = 12'h000;
            11670: color = 12'h000;
            11671: color = 12'h000;
            11672: color = 12'h000;
            11673: color = 12'h000;
            11674: color = 12'h000;
            11675: color = 12'h000;
            11676: color = 12'h000;
            11677: color = 12'h000;
            11678: color = 12'h000;
            11679: color = 12'h000;
            11680: color = 12'h000;
            11681: color = 12'h000;
            11682: color = 12'h000;
            11683: color = 12'h000;
            11684: color = 12'h000;
            11685: color = 12'h000;
            11686: color = 12'h000;
            11687: color = 12'h000;
            11688: color = 12'h000;
            11689: color = 12'h000;
            11690: color = 12'h000;
            11691: color = 12'h000;
            11692: color = 12'h000;
            11693: color = 12'h000;
            11694: color = 12'h000;
            11695: color = 12'h000;
            11696: color = 12'h000;
            11697: color = 12'h000;
            11698: color = 12'h000;
            11699: color = 12'h000;
            11700: color = 12'h000;
            11701: color = 12'h000;
            11702: color = 12'h000;
            11703: color = 12'h000;
            11704: color = 12'h000;
            11705: color = 12'h000;
            11706: color = 12'h000;
            11707: color = 12'h000;
            11708: color = 12'h000;
            11709: color = 12'h000;
            11710: color = 12'h000;
            11711: color = 12'h000;
            11712: color = 12'h000;
            11713: color = 12'h000;
            11714: color = 12'h000;
            11715: color = 12'h000;
            11716: color = 12'h000;
            11717: color = 12'h000;
            11718: color = 12'h000;
            11719: color = 12'h000;
            11720: color = 12'h000;
            11721: color = 12'h000;
            11722: color = 12'h000;
            11723: color = 12'h000;
            11724: color = 12'h000;
            11725: color = 12'h000;
            11726: color = 12'h000;
            11727: color = 12'h000;
            11728: color = 12'h000;
            11729: color = 12'h000;
            11730: color = 12'h000;
            11731: color = 12'h000;
            11732: color = 12'h000;
            11733: color = 12'h000;
            11734: color = 12'h000;
            11735: color = 12'h000;
            11736: color = 12'h000;
            11737: color = 12'h000;
            11738: color = 12'h000;
            11739: color = 12'h000;
            11740: color = 12'h000;
            11741: color = 12'h000;
            11742: color = 12'h000;
            11743: color = 12'h000;
            11744: color = 12'h000;
            11745: color = 12'h000;
            11746: color = 12'h000;
            11747: color = 12'h000;
            11748: color = 12'h000;
            11749: color = 12'h000;
            11750: color = 12'h000;
            11751: color = 12'h000;
            11752: color = 12'h000;
            11753: color = 12'h000;
            11754: color = 12'h000;
            11755: color = 12'h000;
            11756: color = 12'h000;
            11757: color = 12'h000;
            11758: color = 12'h000;
            11759: color = 12'h000;
            11760: color = 12'h000;
            11761: color = 12'h000;
            11762: color = 12'h000;
            11763: color = 12'h000;
            11764: color = 12'h000;
            11765: color = 12'h000;
            11766: color = 12'h000;
            11767: color = 12'h000;
            11768: color = 12'h000;
            11769: color = 12'h000;
            11770: color = 12'h000;
            11771: color = 12'h000;
            11772: color = 12'h000;
            11773: color = 12'h000;
            11774: color = 12'h000;
            11775: color = 12'h000;
            11776: color = 12'h000;
            11777: color = 12'h000;
            11778: color = 12'h000;
            11779: color = 12'h000;
            11780: color = 12'h000;
            11781: color = 12'h000;
            11782: color = 12'h000;
            11783: color = 12'h000;
            11784: color = 12'h000;
            11785: color = 12'h000;
            11786: color = 12'h000;
            11787: color = 12'h000;
            11788: color = 12'h000;
            11789: color = 12'h000;
            11790: color = 12'h000;
            11791: color = 12'h000;
            11792: color = 12'h000;
            11793: color = 12'h000;
            11794: color = 12'h000;
            11795: color = 12'h000;
            11796: color = 12'h000;
            11797: color = 12'h000;
            11798: color = 12'h000;
            11799: color = 12'h000;
            11800: color = 12'h000;
            11801: color = 12'h000;
            11802: color = 12'h000;
            11803: color = 12'h000;
            11804: color = 12'h000;
            11805: color = 12'h000;
            11806: color = 12'h000;
            11807: color = 12'h000;
            11808: color = 12'h000;
            11809: color = 12'h000;
            11810: color = 12'h000;
            11811: color = 12'h000;
            11812: color = 12'h000;
            11813: color = 12'h000;
            11814: color = 12'h000;
            11815: color = 12'h000;
            11816: color = 12'h000;
            11817: color = 12'h000;
            11818: color = 12'h000;
            11819: color = 12'h000;
            11820: color = 12'h000;
            11821: color = 12'h000;
            11822: color = 12'h000;
            11823: color = 12'h000;
            11824: color = 12'h000;
            11825: color = 12'h000;
            11826: color = 12'h000;
            11827: color = 12'h000;
            11828: color = 12'h000;
            11829: color = 12'h000;
            11830: color = 12'h000;
            11831: color = 12'h000;
            11832: color = 12'h000;
            11833: color = 12'h000;
            11834: color = 12'h000;
            11835: color = 12'h000;
            11836: color = 12'h000;
            11837: color = 12'h000;
            11838: color = 12'h000;
            11839: color = 12'h000;
            11840: color = 12'h000;
            11841: color = 12'h000;
            11842: color = 12'h000;
            11843: color = 12'h000;
            11844: color = 12'h000;
            11845: color = 12'h000;
            11846: color = 12'h000;
            11847: color = 12'h000;
            11848: color = 12'h000;
            11849: color = 12'h000;
            11850: color = 12'h000;
            11851: color = 12'h000;
            11852: color = 12'h000;
            11853: color = 12'h000;
            11854: color = 12'h000;
            11855: color = 12'h000;
            11856: color = 12'h000;
            11857: color = 12'h000;
            11858: color = 12'h000;
            11859: color = 12'h000;
            11860: color = 12'h000;
            11861: color = 12'h000;
            11862: color = 12'h000;
            11863: color = 12'h000;
            11864: color = 12'h000;
            11865: color = 12'h000;
            11866: color = 12'h000;
            11867: color = 12'h000;
            11868: color = 12'h000;
            11869: color = 12'h000;
            11870: color = 12'h000;
            11871: color = 12'h000;
            11872: color = 12'h000;
            11873: color = 12'h000;
            11874: color = 12'h000;
            11875: color = 12'h000;
            11876: color = 12'h000;
            11877: color = 12'h000;
            11878: color = 12'h000;
            11879: color = 12'h000;
            11880: color = 12'h000;
            11881: color = 12'h000;
            11882: color = 12'h000;
            11883: color = 12'h000;
            11884: color = 12'h000;
            11885: color = 12'h000;
            11886: color = 12'h000;
            11887: color = 12'h000;
            11888: color = 12'h000;
            11889: color = 12'h000;
            11890: color = 12'h000;
            11891: color = 12'h000;
            11892: color = 12'h000;
            11893: color = 12'h000;
            11894: color = 12'h000;
            11895: color = 12'h000;
            11896: color = 12'h000;
            11897: color = 12'h000;
            11898: color = 12'h000;
            11899: color = 12'h000;
            11900: color = 12'h000;
            11901: color = 12'h000;
            11902: color = 12'h000;
            11903: color = 12'h000;
            11904: color = 12'h000;
            11905: color = 12'h000;
            11906: color = 12'h000;
            11907: color = 12'h000;
            11908: color = 12'h000;
            11909: color = 12'h000;
            11910: color = 12'h000;
            11911: color = 12'h000;
            11912: color = 12'h000;
            11913: color = 12'h000;
            11914: color = 12'h000;
            11915: color = 12'h000;
            11916: color = 12'h000;
            11917: color = 12'h000;
            11918: color = 12'h000;
            11919: color = 12'h000;
            11920: color = 12'h000;
            11921: color = 12'h000;
            11922: color = 12'h000;
            11923: color = 12'h000;
            11924: color = 12'h000;
            11925: color = 12'h000;
            11926: color = 12'h000;
            11927: color = 12'h000;
            11928: color = 12'h000;
            11929: color = 12'h000;
            11930: color = 12'h000;
            11931: color = 12'h000;
            11932: color = 12'h000;
            11933: color = 12'h000;
            11934: color = 12'h000;
            11935: color = 12'h000;
            11936: color = 12'h000;
            11937: color = 12'h000;
            11938: color = 12'h000;
            11939: color = 12'h000;
            11940: color = 12'h000;
            11941: color = 12'h000;
            11942: color = 12'h000;
            11943: color = 12'h000;
            11944: color = 12'h000;
            11945: color = 12'h000;
            11946: color = 12'h000;
            11947: color = 12'h000;
            11948: color = 12'h000;
            11949: color = 12'h000;
            11950: color = 12'h000;
            11951: color = 12'h000;
            11952: color = 12'h000;
            11953: color = 12'h000;
            11954: color = 12'h000;
            11955: color = 12'h000;
            11956: color = 12'h000;
            11957: color = 12'h000;
            11958: color = 12'h000;
            11959: color = 12'h000;
            11960: color = 12'h000;
            11961: color = 12'h000;
            11962: color = 12'h000;
            11963: color = 12'h000;
            11964: color = 12'h000;
            11965: color = 12'h000;
            11966: color = 12'h000;
            11967: color = 12'h000;
            11968: color = 12'h000;
            11969: color = 12'h000;
            11970: color = 12'h000;
            11971: color = 12'h000;
            11972: color = 12'h000;
            11973: color = 12'h000;
            11974: color = 12'h000;
            11975: color = 12'h000;
            11976: color = 12'h000;
            11977: color = 12'h000;
            11978: color = 12'h000;
            11979: color = 12'h000;
            11980: color = 12'h000;
            11981: color = 12'h000;
            11982: color = 12'h000;
            11983: color = 12'h000;
            11984: color = 12'h000;
            11985: color = 12'h000;
            11986: color = 12'h000;
            11987: color = 12'h000;
            11988: color = 12'h000;
            11989: color = 12'h000;
            11990: color = 12'h000;
            11991: color = 12'h000;
            11992: color = 12'h000;
            11993: color = 12'h000;
            11994: color = 12'h000;
            11995: color = 12'h000;
            11996: color = 12'h000;
            11997: color = 12'h000;
            11998: color = 12'h000;
            11999: color = 12'h000;
            12000: color = 12'h000;
            12001: color = 12'h000;
            12002: color = 12'h000;
            12003: color = 12'h000;
            12004: color = 12'h000;
            12005: color = 12'h000;
            12006: color = 12'h000;
            12007: color = 12'h000;
            12008: color = 12'h000;
            12009: color = 12'h000;
            12010: color = 12'h000;
            12011: color = 12'h000;
            12012: color = 12'h000;
            12013: color = 12'h000;
            12014: color = 12'h000;
            12015: color = 12'h000;
            12016: color = 12'h000;
            12017: color = 12'h000;
            12018: color = 12'h000;
            12019: color = 12'h000;
            12020: color = 12'h000;
            12021: color = 12'h000;
            12022: color = 12'h000;
            12023: color = 12'h000;
            12024: color = 12'h000;
            12025: color = 12'h000;
            12026: color = 12'h000;
            12027: color = 12'h000;
            12028: color = 12'h000;
            12029: color = 12'h000;
            12030: color = 12'h000;
            12031: color = 12'h000;
            12032: color = 12'h000;
            12033: color = 12'h000;
            12034: color = 12'h000;
            12035: color = 12'h000;
            12036: color = 12'h000;
            12037: color = 12'h000;
            12038: color = 12'h000;
            12039: color = 12'h000;
            12040: color = 12'h000;
            12041: color = 12'h000;
            12042: color = 12'h000;
            12043: color = 12'h000;
            12044: color = 12'h000;
            12045: color = 12'h000;
            12046: color = 12'h000;
            12047: color = 12'h000;
            12048: color = 12'h000;
            12049: color = 12'h000;
            12050: color = 12'h000;
            12051: color = 12'h000;
            12052: color = 12'h000;
            12053: color = 12'h000;
            12054: color = 12'h000;
            12055: color = 12'h000;
            12056: color = 12'h000;
            12057: color = 12'h000;
            12058: color = 12'h000;
            12059: color = 12'h000;
            12060: color = 12'h000;
            12061: color = 12'h000;
            12062: color = 12'h000;
            12063: color = 12'h000;
            12064: color = 12'h000;
            12065: color = 12'h000;
            12066: color = 12'h000;
            12067: color = 12'h000;
            12068: color = 12'h000;
            12069: color = 12'h000;
            12070: color = 12'h000;
            12071: color = 12'h000;
            12072: color = 12'h000;
            12073: color = 12'h000;
            12074: color = 12'h000;
            12075: color = 12'h000;
            12076: color = 12'h000;
            12077: color = 12'h000;
            12078: color = 12'h000;
            12079: color = 12'h000;
            12080: color = 12'h000;
            12081: color = 12'h000;
            12082: color = 12'h000;
            12083: color = 12'h000;
            12084: color = 12'h000;
            12085: color = 12'h000;
            12086: color = 12'h000;
            12087: color = 12'h000;
            12088: color = 12'h000;
            12089: color = 12'h000;
            12090: color = 12'h000;
            12091: color = 12'h000;
            12092: color = 12'h000;
            12093: color = 12'h000;
            12094: color = 12'h000;
            12095: color = 12'h000;
            12096: color = 12'h000;
            12097: color = 12'h000;
            12098: color = 12'h000;
            12099: color = 12'h000;
            12100: color = 12'h000;
            12101: color = 12'h000;
            12102: color = 12'h000;
            12103: color = 12'h000;
            12104: color = 12'h000;
            12105: color = 12'h000;
            12106: color = 12'h000;
            12107: color = 12'h000;
            12108: color = 12'h000;
            12109: color = 12'h000;
            12110: color = 12'h000;
            12111: color = 12'h000;
            12112: color = 12'h000;
            12113: color = 12'h000;
            12114: color = 12'h000;
            12115: color = 12'h000;
            12116: color = 12'h000;
            12117: color = 12'h000;
            12118: color = 12'h000;
            12119: color = 12'h000;
            12120: color = 12'h000;
            12121: color = 12'h000;
            12122: color = 12'h000;
            12123: color = 12'h000;
            12124: color = 12'h000;
            12125: color = 12'h000;
            12126: color = 12'h000;
            12127: color = 12'h000;
            12128: color = 12'h000;
            12129: color = 12'h000;
            12130: color = 12'h000;
            12131: color = 12'h000;
            12132: color = 12'h000;
            12133: color = 12'h000;
            12134: color = 12'h000;
            12135: color = 12'h000;
            12136: color = 12'h000;
            12137: color = 12'h000;
            12138: color = 12'h000;
            12139: color = 12'h000;
            12140: color = 12'h000;
            12141: color = 12'h000;
            12142: color = 12'h000;
            12143: color = 12'h000;
            12144: color = 12'h000;
            12145: color = 12'h000;
            12146: color = 12'h000;
            12147: color = 12'h000;
            12148: color = 12'h000;
            12149: color = 12'h000;
            12150: color = 12'h000;
            12151: color = 12'h000;
            12152: color = 12'h000;
            12153: color = 12'h000;
            12154: color = 12'h000;
            12155: color = 12'h000;
            12156: color = 12'h000;
            12157: color = 12'h000;
            12158: color = 12'h000;
            12159: color = 12'h000;
            12160: color = 12'h000;
            12161: color = 12'h000;
            12162: color = 12'h000;
            12163: color = 12'h000;
            12164: color = 12'h000;
            12165: color = 12'h000;
            12166: color = 12'h000;
            12167: color = 12'h000;
            12168: color = 12'h000;
            12169: color = 12'h000;
            12170: color = 12'h000;
            12171: color = 12'h000;
            12172: color = 12'h000;
            12173: color = 12'h000;
            12174: color = 12'h000;
            12175: color = 12'h000;
            12176: color = 12'h000;
            12177: color = 12'h000;
            12178: color = 12'h000;
            12179: color = 12'h000;
            12180: color = 12'h000;
            12181: color = 12'h000;
            12182: color = 12'h000;
            12183: color = 12'h000;
            12184: color = 12'h000;
            12185: color = 12'h000;
            12186: color = 12'h000;
            12187: color = 12'h000;
            12188: color = 12'h000;
            12189: color = 12'h000;
            12190: color = 12'h000;
            12191: color = 12'h000;
            12192: color = 12'h000;
            12193: color = 12'h000;
            12194: color = 12'h000;
            12195: color = 12'h000;
            12196: color = 12'h000;
            12197: color = 12'h000;
            12198: color = 12'h000;
            12199: color = 12'h000;
            12200: color = 12'h000;
            12201: color = 12'h000;
            12202: color = 12'h000;
            12203: color = 12'h000;
            12204: color = 12'h000;
            12205: color = 12'h000;
            12206: color = 12'h000;
            12207: color = 12'h000;
            12208: color = 12'h000;
            12209: color = 12'h000;
            12210: color = 12'h000;
            12211: color = 12'h000;
            12212: color = 12'h000;
            12213: color = 12'h000;
            12214: color = 12'h000;
            12215: color = 12'h000;
            12216: color = 12'h000;
            12217: color = 12'h000;
            12218: color = 12'h000;
            12219: color = 12'h000;
            12220: color = 12'h000;
            12221: color = 12'h000;
            12222: color = 12'h000;
            12223: color = 12'h000;
            12224: color = 12'h000;
            12225: color = 12'h000;
            12226: color = 12'h000;
            12227: color = 12'h000;
            12228: color = 12'h000;
            12229: color = 12'h000;
            12230: color = 12'h000;
            12231: color = 12'h000;
            12232: color = 12'h000;
            12233: color = 12'h000;
            12234: color = 12'h000;
            12235: color = 12'h000;
            12236: color = 12'h000;
            12237: color = 12'h000;
            12238: color = 12'h000;
            12239: color = 12'h000;
            12240: color = 12'h000;
            12241: color = 12'h000;
            12242: color = 12'h000;
            12243: color = 12'h000;
            12244: color = 12'h000;
            12245: color = 12'h000;
            12246: color = 12'h000;
            12247: color = 12'h000;
            12248: color = 12'h000;
            12249: color = 12'h000;
            12250: color = 12'h000;
            12251: color = 12'h000;
            12252: color = 12'h000;
            12253: color = 12'h000;
            12254: color = 12'h000;
            12255: color = 12'h000;
            12256: color = 12'h000;
            12257: color = 12'h000;
            12258: color = 12'h000;
            12259: color = 12'h000;
            12260: color = 12'h000;
            12261: color = 12'h000;
            12262: color = 12'h000;
            12263: color = 12'h000;
            12264: color = 12'h000;
            12265: color = 12'h000;
            12266: color = 12'h000;
            12267: color = 12'h000;
            12268: color = 12'h000;
            12269: color = 12'h000;
            12270: color = 12'h000;
            12271: color = 12'h000;
            12272: color = 12'h000;
            12273: color = 12'h000;
            12274: color = 12'h000;
            12275: color = 12'h000;
            12276: color = 12'h000;
            12277: color = 12'h000;
            12278: color = 12'h000;
            12279: color = 12'h000;
            12280: color = 12'h000;
            12281: color = 12'h000;
            12282: color = 12'h000;
            12283: color = 12'h000;
            12284: color = 12'h000;
            12285: color = 12'h000;
            12286: color = 12'h000;
            12287: color = 12'h000;
            12288: color = 12'h000;
            12289: color = 12'h000;
            12290: color = 12'h000;
            12291: color = 12'h000;
            12292: color = 12'h000;
            12293: color = 12'h000;
            12294: color = 12'h000;
            12295: color = 12'h000;
            12296: color = 12'h000;
            12297: color = 12'h000;
            12298: color = 12'h000;
            12299: color = 12'h000;
            12300: color = 12'h000;
            12301: color = 12'h000;
            12302: color = 12'h000;
            12303: color = 12'h000;
            12304: color = 12'h000;
            12305: color = 12'h000;
            12306: color = 12'h000;
            12307: color = 12'h000;
            12308: color = 12'h000;
            12309: color = 12'h000;
            12310: color = 12'h000;
            12311: color = 12'h000;
            12312: color = 12'h000;
            12313: color = 12'h000;
            12314: color = 12'h000;
            12315: color = 12'h000;
            12316: color = 12'h000;
            12317: color = 12'h000;
            12318: color = 12'h000;
            12319: color = 12'h000;
            12320: color = 12'h000;
            12321: color = 12'h000;
            12322: color = 12'h000;
            12323: color = 12'h000;
            12324: color = 12'h000;
            12325: color = 12'h000;
            12326: color = 12'h000;
            12327: color = 12'h000;
            12328: color = 12'h000;
            12329: color = 12'h000;
            12330: color = 12'h000;
            12331: color = 12'h000;
            12332: color = 12'h000;
            12333: color = 12'h000;
            12334: color = 12'h000;
            12335: color = 12'h000;
            12336: color = 12'h000;
            12337: color = 12'h000;
            12338: color = 12'h000;
            12339: color = 12'h000;
            12340: color = 12'h000;
            12341: color = 12'h000;
            12342: color = 12'h000;
            12343: color = 12'h000;
            12344: color = 12'h000;
            12345: color = 12'h000;
            12346: color = 12'h000;
            12347: color = 12'h000;
            12348: color = 12'h000;
            12349: color = 12'h000;
            12350: color = 12'h000;
            12351: color = 12'h000;
            12352: color = 12'h000;
            12353: color = 12'h000;
            12354: color = 12'h000;
            12355: color = 12'h000;
            12356: color = 12'h000;
            12357: color = 12'h000;
            12358: color = 12'h000;
            12359: color = 12'h000;
            12360: color = 12'h000;
            12361: color = 12'h000;
            12362: color = 12'h000;
            12363: color = 12'h000;
            12364: color = 12'h000;
            12365: color = 12'h000;
            12366: color = 12'h000;
            12367: color = 12'h000;
            12368: color = 12'h000;
            12369: color = 12'h000;
            12370: color = 12'h000;
            12371: color = 12'h000;
            12372: color = 12'h000;
            12373: color = 12'h000;
            12374: color = 12'h000;
            12375: color = 12'h000;
            12376: color = 12'h000;
            12377: color = 12'h000;
            12378: color = 12'h000;
            12379: color = 12'h000;
            12380: color = 12'h000;
            12381: color = 12'h000;
            12382: color = 12'h000;
            12383: color = 12'h000;
            12384: color = 12'h000;
            12385: color = 12'h000;
            12386: color = 12'h000;
            12387: color = 12'h000;
            12388: color = 12'h000;
            12389: color = 12'h000;
            12390: color = 12'h000;
            12391: color = 12'h000;
            12392: color = 12'h000;
            12393: color = 12'h000;
            12394: color = 12'h000;
            12395: color = 12'h000;
            12396: color = 12'h000;
            12397: color = 12'h000;
            12398: color = 12'h000;
            12399: color = 12'h000;
            12400: color = 12'h000;
            12401: color = 12'h000;
            12402: color = 12'h000;
            12403: color = 12'h000;
            12404: color = 12'h000;
            12405: color = 12'h000;
            12406: color = 12'h000;
            12407: color = 12'h000;
            12408: color = 12'h000;
            12409: color = 12'h000;
            12410: color = 12'h000;
            12411: color = 12'h000;
            12412: color = 12'h000;
            12413: color = 12'h000;
            12414: color = 12'h000;
            12415: color = 12'h000;
            12416: color = 12'h000;
            12417: color = 12'h000;
            12418: color = 12'h000;
            12419: color = 12'h000;
            12420: color = 12'h000;
            12421: color = 12'h000;
            12422: color = 12'h000;
            12423: color = 12'h000;
            12424: color = 12'h000;
            12425: color = 12'h000;
            12426: color = 12'h000;
            12427: color = 12'h000;
            12428: color = 12'h000;
            12429: color = 12'h000;
            12430: color = 12'h000;
            12431: color = 12'h000;
            12432: color = 12'h000;
            12433: color = 12'h000;
            12434: color = 12'h000;
            12435: color = 12'h000;
            12436: color = 12'h000;
            12437: color = 12'h000;
            12438: color = 12'h000;
            12439: color = 12'h000;
            12440: color = 12'h000;
            12441: color = 12'h000;
            12442: color = 12'h000;
            12443: color = 12'h000;
            12444: color = 12'h000;
            12445: color = 12'h000;
            12446: color = 12'h000;
            12447: color = 12'h000;
            12448: color = 12'h000;
            12449: color = 12'h000;
            12450: color = 12'h000;
            12451: color = 12'h000;
            12452: color = 12'h000;
            12453: color = 12'h000;
            12454: color = 12'h000;
            12455: color = 12'h000;
            12456: color = 12'h000;
            12457: color = 12'h000;
            12458: color = 12'h000;
            12459: color = 12'h000;
            12460: color = 12'h000;
            12461: color = 12'h000;
            12462: color = 12'h000;
            12463: color = 12'h000;
            12464: color = 12'h000;
            12465: color = 12'h000;
            12466: color = 12'h000;
            12467: color = 12'h000;
            12468: color = 12'h000;
            12469: color = 12'h000;
            12470: color = 12'h000;
            12471: color = 12'h000;
            12472: color = 12'h000;
            12473: color = 12'h000;
            12474: color = 12'h000;
            12475: color = 12'h000;
            12476: color = 12'h000;
            12477: color = 12'h000;
            12478: color = 12'h000;
            12479: color = 12'h000;
            12480: color = 12'h000;
            12481: color = 12'h000;
            12482: color = 12'h000;
            12483: color = 12'h000;
            12484: color = 12'h000;
            12485: color = 12'h000;
            12486: color = 12'h000;
            12487: color = 12'h000;
            12488: color = 12'h000;
            12489: color = 12'h000;
            12490: color = 12'h000;
            12491: color = 12'h000;
            12492: color = 12'h000;
            12493: color = 12'h000;
            12494: color = 12'h000;
            12495: color = 12'h000;
            12496: color = 12'h000;
            12497: color = 12'h000;
            12498: color = 12'h000;
            12499: color = 12'h000;
            12500: color = 12'h000;
            12501: color = 12'h000;
            12502: color = 12'h000;
            12503: color = 12'h000;
            12504: color = 12'h000;
            12505: color = 12'h000;
            12506: color = 12'h000;
            12507: color = 12'h000;
            12508: color = 12'h000;
            12509: color = 12'h000;
            12510: color = 12'h000;
            12511: color = 12'h000;
            12512: color = 12'h000;
            12513: color = 12'h000;
            12514: color = 12'h000;
            12515: color = 12'h000;
            12516: color = 12'h000;
            12517: color = 12'h000;
            12518: color = 12'h000;
            12519: color = 12'h000;
            12520: color = 12'h000;
            12521: color = 12'h000;
            12522: color = 12'h000;
            12523: color = 12'h000;
            12524: color = 12'h000;
            12525: color = 12'h000;
            12526: color = 12'h000;
            12527: color = 12'h000;
            12528: color = 12'h000;
            12529: color = 12'h000;
            12530: color = 12'h000;
            12531: color = 12'h000;
            12532: color = 12'h000;
            12533: color = 12'h000;
            12534: color = 12'h000;
            12535: color = 12'h000;
            12536: color = 12'h000;
            12537: color = 12'h000;
            12538: color = 12'h000;
            12539: color = 12'h000;
            12540: color = 12'h000;
            12541: color = 12'h000;
            12542: color = 12'h000;
            12543: color = 12'h000;
            12544: color = 12'h000;
            12545: color = 12'h000;
            12546: color = 12'h000;
            12547: color = 12'h000;
            12548: color = 12'h000;
            12549: color = 12'h000;
            12550: color = 12'h000;
            12551: color = 12'h000;
            12552: color = 12'h000;
            12553: color = 12'h000;
            12554: color = 12'h000;
            12555: color = 12'h000;
            12556: color = 12'h000;
            12557: color = 12'h000;
            12558: color = 12'h000;
            12559: color = 12'h000;
            12560: color = 12'h000;
            12561: color = 12'h000;
            12562: color = 12'h000;
            12563: color = 12'h000;
            12564: color = 12'h000;
            12565: color = 12'h000;
            12566: color = 12'h000;
            12567: color = 12'h000;
            12568: color = 12'h000;
            12569: color = 12'h000;
            12570: color = 12'h000;
            12571: color = 12'h000;
            12572: color = 12'h000;
            12573: color = 12'h000;
            12574: color = 12'h000;
            12575: color = 12'h000;
            12576: color = 12'h000;
            12577: color = 12'h000;
            12578: color = 12'h000;
            12579: color = 12'h000;
            12580: color = 12'h000;
            12581: color = 12'h000;
            12582: color = 12'h000;
            12583: color = 12'h000;
            12584: color = 12'h000;
            12585: color = 12'h000;
            12586: color = 12'h000;
            12587: color = 12'h000;
            12588: color = 12'h000;
            12589: color = 12'h000;
            12590: color = 12'h000;
            12591: color = 12'h000;
            12592: color = 12'h000;
            12593: color = 12'h000;
            12594: color = 12'h000;
            12595: color = 12'h000;
            12596: color = 12'h000;
            12597: color = 12'h000;
            12598: color = 12'h000;
            12599: color = 12'h000;
            12600: color = 12'h000;
            12601: color = 12'h000;
            12602: color = 12'h000;
            12603: color = 12'h000;
            12604: color = 12'h000;
            12605: color = 12'h000;
            12606: color = 12'h000;
            12607: color = 12'h000;
            12608: color = 12'h000;
            12609: color = 12'h000;
            12610: color = 12'h000;
            12611: color = 12'h000;
            12612: color = 12'h000;
            12613: color = 12'h000;
            12614: color = 12'h000;
            12615: color = 12'h000;
            12616: color = 12'h000;
            12617: color = 12'h000;
            12618: color = 12'h000;
            12619: color = 12'h000;
            12620: color = 12'h000;
            12621: color = 12'h000;
            12622: color = 12'h000;
            12623: color = 12'h000;
            12624: color = 12'h000;
            12625: color = 12'h000;
            12626: color = 12'h000;
            12627: color = 12'h000;
            12628: color = 12'h000;
            12629: color = 12'h000;
            12630: color = 12'h000;
            12631: color = 12'h000;
            12632: color = 12'h000;
            12633: color = 12'h000;
            12634: color = 12'h000;
            12635: color = 12'h000;
            12636: color = 12'h000;
            12637: color = 12'h000;
            12638: color = 12'h000;
            12639: color = 12'h000;
            12640: color = 12'h000;
            12641: color = 12'h000;
            12642: color = 12'h000;
            12643: color = 12'h000;
            12644: color = 12'h000;
            12645: color = 12'h000;
            12646: color = 12'h000;
            12647: color = 12'h000;
            12648: color = 12'h000;
            12649: color = 12'h000;
            12650: color = 12'h000;
            12651: color = 12'h000;
            12652: color = 12'h000;
            12653: color = 12'h000;
            12654: color = 12'h000;
            12655: color = 12'h000;
            12656: color = 12'h000;
            12657: color = 12'h000;
            12658: color = 12'h000;
            12659: color = 12'h000;
            12660: color = 12'h000;
            12661: color = 12'h000;
            12662: color = 12'h000;
            12663: color = 12'h000;
            12664: color = 12'h000;
            12665: color = 12'h000;
            12666: color = 12'h000;
            12667: color = 12'h000;
            12668: color = 12'h000;
            12669: color = 12'h000;
            12670: color = 12'h000;
            12671: color = 12'h000;
            12672: color = 12'h000;
            12673: color = 12'h000;
            12674: color = 12'h000;
            12675: color = 12'h000;
            12676: color = 12'h000;
            12677: color = 12'h000;
            12678: color = 12'h000;
            12679: color = 12'h000;
            12680: color = 12'h000;
            12681: color = 12'h000;
            12682: color = 12'h000;
            12683: color = 12'h000;
            12684: color = 12'h000;
            12685: color = 12'h000;
            12686: color = 12'h000;
            12687: color = 12'h000;
            12688: color = 12'h000;
            12689: color = 12'h000;
            12690: color = 12'h000;
            12691: color = 12'h000;
            12692: color = 12'h000;
            12693: color = 12'h000;
            12694: color = 12'h000;
            12695: color = 12'h000;
            12696: color = 12'h000;
            12697: color = 12'h000;
            12698: color = 12'h000;
            12699: color = 12'h000;
            12700: color = 12'h000;
            12701: color = 12'h000;
            12702: color = 12'h000;
            12703: color = 12'h000;
            12704: color = 12'h000;
            12705: color = 12'h000;
            12706: color = 12'h000;
            12707: color = 12'h000;
            12708: color = 12'h000;
            12709: color = 12'h000;
            12710: color = 12'h000;
            12711: color = 12'h000;
            12712: color = 12'h000;
            12713: color = 12'h000;
            12714: color = 12'h000;
            12715: color = 12'h000;
            12716: color = 12'h000;
            12717: color = 12'h000;
            12718: color = 12'h000;
            12719: color = 12'h000;
            12720: color = 12'h000;
            12721: color = 12'h000;
            12722: color = 12'h000;
            12723: color = 12'h000;
            12724: color = 12'h000;
            12725: color = 12'h000;
            12726: color = 12'h000;
            12727: color = 12'h000;
            12728: color = 12'h000;
            12729: color = 12'h000;
            12730: color = 12'h000;
            12731: color = 12'h000;
            12732: color = 12'h000;
            12733: color = 12'h000;
            12734: color = 12'h000;
            12735: color = 12'h000;
            12736: color = 12'h000;
            12737: color = 12'h000;
            12738: color = 12'h000;
            12739: color = 12'h000;
            12740: color = 12'h000;
            12741: color = 12'h000;
            12742: color = 12'h000;
            12743: color = 12'h000;
            12744: color = 12'h000;
            12745: color = 12'h000;
            12746: color = 12'h000;
            12747: color = 12'h000;
            12748: color = 12'h000;
            12749: color = 12'h000;
            12750: color = 12'h000;
            12751: color = 12'h000;
            12752: color = 12'h000;
            12753: color = 12'h000;
            12754: color = 12'h000;
            12755: color = 12'h000;
            12756: color = 12'h000;
            12757: color = 12'h000;
            12758: color = 12'h000;
            12759: color = 12'h000;
            12760: color = 12'h000;
            12761: color = 12'h000;
            12762: color = 12'h000;
            12763: color = 12'h000;
            12764: color = 12'h000;
            12765: color = 12'h000;
            12766: color = 12'h000;
            12767: color = 12'h000;
            12768: color = 12'h000;
            12769: color = 12'h000;
            12770: color = 12'h000;
            12771: color = 12'h000;
            12772: color = 12'h000;
            12773: color = 12'h000;
            12774: color = 12'h000;
            12775: color = 12'h000;
            12776: color = 12'h000;
            12777: color = 12'h000;
            12778: color = 12'h000;
            12779: color = 12'h000;
            12780: color = 12'h000;
            12781: color = 12'h000;
            12782: color = 12'h000;
            12783: color = 12'h000;
            12784: color = 12'h000;
            12785: color = 12'h000;
            12786: color = 12'h000;
            12787: color = 12'h000;
            12788: color = 12'h000;
            12789: color = 12'h000;
            12790: color = 12'h000;
            12791: color = 12'h000;
            12792: color = 12'h000;
            12793: color = 12'h000;
            12794: color = 12'h000;
            12795: color = 12'h000;
            12796: color = 12'h000;
            12797: color = 12'h000;
            12798: color = 12'h000;
            12799: color = 12'h000;
            12800: color = 12'h000;
            12801: color = 12'h000;
            12802: color = 12'h000;
            12803: color = 12'h000;
            12804: color = 12'h000;
            12805: color = 12'h000;
            12806: color = 12'h000;
            12807: color = 12'h000;
            12808: color = 12'h000;
            12809: color = 12'h000;
            12810: color = 12'h000;
            12811: color = 12'h000;
            12812: color = 12'h000;
            12813: color = 12'h000;
            12814: color = 12'h000;
            12815: color = 12'h000;
            12816: color = 12'h000;
            12817: color = 12'h000;
            12818: color = 12'h000;
            12819: color = 12'h000;
            12820: color = 12'h000;
            12821: color = 12'h000;
            12822: color = 12'h000;
            12823: color = 12'h000;
            12824: color = 12'h000;
            12825: color = 12'h000;
            12826: color = 12'h000;
            12827: color = 12'h000;
            12828: color = 12'h000;
            12829: color = 12'h000;
            12830: color = 12'h000;
            12831: color = 12'h000;
            12832: color = 12'h000;
            12833: color = 12'h000;
            12834: color = 12'h000;
            12835: color = 12'h000;
            12836: color = 12'h000;
            12837: color = 12'h000;
            12838: color = 12'h000;
            12839: color = 12'h000;
            12840: color = 12'h000;
            12841: color = 12'h000;
            12842: color = 12'h000;
            12843: color = 12'h000;
            12844: color = 12'h000;
            12845: color = 12'h000;
            12846: color = 12'h000;
            12847: color = 12'h000;
            12848: color = 12'h000;
            12849: color = 12'h000;
            12850: color = 12'h000;
            12851: color = 12'h000;
            12852: color = 12'h000;
            12853: color = 12'h000;
            12854: color = 12'h000;
            12855: color = 12'h000;
            12856: color = 12'h000;
            12857: color = 12'h000;
            12858: color = 12'h000;
            12859: color = 12'h000;
            12860: color = 12'h000;
            12861: color = 12'h000;
            12862: color = 12'h000;
            12863: color = 12'h000;
            12864: color = 12'h000;
            12865: color = 12'h000;
            12866: color = 12'h000;
            12867: color = 12'h000;
            12868: color = 12'h000;
            12869: color = 12'h000;
            12870: color = 12'h000;
            12871: color = 12'h000;
            12872: color = 12'h000;
            12873: color = 12'h000;
            12874: color = 12'h000;
            12875: color = 12'h000;
            12876: color = 12'h000;
            12877: color = 12'h000;
            12878: color = 12'h000;
            12879: color = 12'h000;
            12880: color = 12'h000;
            12881: color = 12'h000;
            12882: color = 12'h000;
            12883: color = 12'h000;
            12884: color = 12'h000;
            12885: color = 12'h000;
            12886: color = 12'h000;
            12887: color = 12'h000;
            12888: color = 12'h000;
            12889: color = 12'h000;
            12890: color = 12'h000;
            12891: color = 12'h000;
            12892: color = 12'h000;
            12893: color = 12'h000;
            12894: color = 12'h000;
            12895: color = 12'h000;
            12896: color = 12'h000;
            12897: color = 12'h000;
            12898: color = 12'h000;
            12899: color = 12'h000;
            12900: color = 12'h000;
            12901: color = 12'h000;
            12902: color = 12'h000;
            12903: color = 12'h000;
            12904: color = 12'h000;
            12905: color = 12'h000;
            12906: color = 12'h000;
            12907: color = 12'h000;
            12908: color = 12'h000;
            12909: color = 12'h000;
            12910: color = 12'h000;
            12911: color = 12'h000;
            12912: color = 12'h000;
            12913: color = 12'h000;
            12914: color = 12'h000;
            12915: color = 12'h000;
            12916: color = 12'h000;
            12917: color = 12'h000;
            12918: color = 12'h000;
            12919: color = 12'h000;
            12920: color = 12'h000;
            12921: color = 12'h000;
            12922: color = 12'h000;
            12923: color = 12'h000;
            12924: color = 12'h000;
            12925: color = 12'h000;
            12926: color = 12'h000;
            12927: color = 12'h000;
            12928: color = 12'h000;
            12929: color = 12'h000;
            12930: color = 12'h000;
            12931: color = 12'h000;
            12932: color = 12'h000;
            12933: color = 12'h000;
            12934: color = 12'h000;
            12935: color = 12'h000;
            12936: color = 12'h000;
            12937: color = 12'h000;
            12938: color = 12'h000;
            12939: color = 12'h000;
            12940: color = 12'h000;
            12941: color = 12'h000;
            12942: color = 12'h000;
            12943: color = 12'h000;
            12944: color = 12'h000;
            12945: color = 12'h000;
            12946: color = 12'h000;
            12947: color = 12'h000;
            12948: color = 12'h000;
            12949: color = 12'h000;
            12950: color = 12'h000;
            12951: color = 12'h000;
            12952: color = 12'h000;
            12953: color = 12'h000;
            12954: color = 12'h000;
            12955: color = 12'h000;
            12956: color = 12'h000;
            12957: color = 12'h000;
            12958: color = 12'h000;
            12959: color = 12'h000;
            12960: color = 12'h000;
            12961: color = 12'h000;
            12962: color = 12'h000;
            12963: color = 12'h000;
            12964: color = 12'h000;
            12965: color = 12'h000;
            12966: color = 12'h000;
            12967: color = 12'h000;
            12968: color = 12'h000;
            12969: color = 12'h000;
            12970: color = 12'h000;
            12971: color = 12'h000;
            12972: color = 12'h000;
            12973: color = 12'h000;
            12974: color = 12'h000;
            12975: color = 12'h000;
            12976: color = 12'h000;
            12977: color = 12'h000;
            12978: color = 12'h000;
            12979: color = 12'h000;
            12980: color = 12'h000;
            12981: color = 12'h000;
            12982: color = 12'h000;
            12983: color = 12'h000;
            12984: color = 12'h000;
            12985: color = 12'h000;
            12986: color = 12'h000;
            12987: color = 12'h000;
            12988: color = 12'h000;
            12989: color = 12'h000;
            12990: color = 12'h000;
            12991: color = 12'h000;
            12992: color = 12'h000;
            12993: color = 12'h000;
            12994: color = 12'h000;
            12995: color = 12'h000;
            12996: color = 12'h000;
            12997: color = 12'h000;
            12998: color = 12'h000;
            12999: color = 12'h000;
            13000: color = 12'h000;
            13001: color = 12'h000;
            13002: color = 12'h000;
            13003: color = 12'h000;
            13004: color = 12'h000;
            13005: color = 12'h000;
            13006: color = 12'h000;
            13007: color = 12'h000;
            13008: color = 12'h000;
            13009: color = 12'h000;
            13010: color = 12'h000;
            13011: color = 12'h000;
            13012: color = 12'h000;
            13013: color = 12'h000;
            13014: color = 12'h000;
            13015: color = 12'h000;
            13016: color = 12'h000;
            13017: color = 12'h000;
            13018: color = 12'h000;
            13019: color = 12'h000;
            13020: color = 12'h000;
            13021: color = 12'h000;
            13022: color = 12'h000;
            13023: color = 12'h000;
            13024: color = 12'h000;
            13025: color = 12'h000;
            13026: color = 12'h000;
            13027: color = 12'h000;
            13028: color = 12'h000;
            13029: color = 12'h000;
            13030: color = 12'h000;
            13031: color = 12'h000;
            13032: color = 12'h000;
            13033: color = 12'h000;
            13034: color = 12'h000;
            13035: color = 12'h000;
            13036: color = 12'h000;
            13037: color = 12'h000;
            13038: color = 12'h000;
            13039: color = 12'h000;
            13040: color = 12'h000;
            13041: color = 12'h000;
            13042: color = 12'h000;
            13043: color = 12'h000;
            13044: color = 12'h000;
            13045: color = 12'h000;
            13046: color = 12'h000;
            13047: color = 12'h000;
            13048: color = 12'h000;
            13049: color = 12'h000;
            13050: color = 12'h000;
            13051: color = 12'h000;
            13052: color = 12'h000;
            13053: color = 12'h000;
            13054: color = 12'h000;
            13055: color = 12'h000;
            13056: color = 12'h000;
            13057: color = 12'h000;
            13058: color = 12'h000;
            13059: color = 12'h000;
            13060: color = 12'h000;
            13061: color = 12'h000;
            13062: color = 12'h000;
            13063: color = 12'h000;
            13064: color = 12'h000;
            13065: color = 12'h000;
            13066: color = 12'h000;
            13067: color = 12'h000;
            13068: color = 12'h000;
            13069: color = 12'h000;
            13070: color = 12'h000;
            13071: color = 12'h000;
            13072: color = 12'h000;
            13073: color = 12'h000;
            13074: color = 12'h000;
            13075: color = 12'h000;
            13076: color = 12'h000;
            13077: color = 12'h000;
            13078: color = 12'h000;
            13079: color = 12'h000;
            13080: color = 12'h000;
            13081: color = 12'h000;
            13082: color = 12'h000;
            13083: color = 12'h000;
            13084: color = 12'h000;
            13085: color = 12'h000;
            13086: color = 12'h000;
            13087: color = 12'h000;
            13088: color = 12'h000;
            13089: color = 12'h000;
            13090: color = 12'h000;
            13091: color = 12'h000;
            13092: color = 12'h000;
            13093: color = 12'h000;
            13094: color = 12'h000;
            13095: color = 12'h000;
            13096: color = 12'h000;
            13097: color = 12'h000;
            13098: color = 12'h000;
            13099: color = 12'h000;
            13100: color = 12'h000;
            13101: color = 12'h000;
            13102: color = 12'h000;
            13103: color = 12'h000;
            13104: color = 12'h000;
            13105: color = 12'h000;
            13106: color = 12'h000;
            13107: color = 12'h000;
            13108: color = 12'h000;
            13109: color = 12'h000;
            13110: color = 12'h000;
            13111: color = 12'h000;
            13112: color = 12'h000;
            13113: color = 12'h000;
            13114: color = 12'h000;
            13115: color = 12'h000;
            13116: color = 12'h000;
            13117: color = 12'h000;
            13118: color = 12'h000;
            13119: color = 12'h000;
            13120: color = 12'h000;
            13121: color = 12'h000;
            13122: color = 12'h000;
            13123: color = 12'h000;
            13124: color = 12'h000;
            13125: color = 12'h000;
            13126: color = 12'h000;
            13127: color = 12'h000;
            13128: color = 12'h000;
            13129: color = 12'h000;
            13130: color = 12'h000;
            13131: color = 12'h000;
            13132: color = 12'h000;
            13133: color = 12'h000;
            13134: color = 12'h000;
            13135: color = 12'h000;
            13136: color = 12'h000;
            13137: color = 12'h000;
            13138: color = 12'h000;
            13139: color = 12'h000;
            13140: color = 12'h000;
            13141: color = 12'h000;
            13142: color = 12'h000;
            13143: color = 12'h000;
            13144: color = 12'h000;
            13145: color = 12'h000;
            13146: color = 12'h000;
            13147: color = 12'h000;
            13148: color = 12'h000;
            13149: color = 12'h000;
            13150: color = 12'h000;
            13151: color = 12'h000;
            13152: color = 12'h000;
            13153: color = 12'h000;
            13154: color = 12'h000;
            13155: color = 12'h000;
            13156: color = 12'h000;
            13157: color = 12'h000;
            13158: color = 12'h000;
            13159: color = 12'h000;
            13160: color = 12'h000;
            13161: color = 12'h000;
            13162: color = 12'h000;
            13163: color = 12'h000;
            13164: color = 12'h000;
            13165: color = 12'h000;
            13166: color = 12'h000;
            13167: color = 12'h000;
            13168: color = 12'h000;
            13169: color = 12'h000;
            13170: color = 12'h000;
            13171: color = 12'h000;
            13172: color = 12'h000;
            13173: color = 12'h000;
            13174: color = 12'h000;
            13175: color = 12'h000;
            13176: color = 12'h000;
            13177: color = 12'h000;
            13178: color = 12'h000;
            13179: color = 12'h000;
            13180: color = 12'h000;
            13181: color = 12'h000;
            13182: color = 12'h000;
            13183: color = 12'h000;
            13184: color = 12'h000;
            13185: color = 12'h000;
            13186: color = 12'h000;
            13187: color = 12'h000;
            13188: color = 12'h000;
            13189: color = 12'h000;
            13190: color = 12'h000;
            13191: color = 12'h000;
            13192: color = 12'h000;
            13193: color = 12'h000;
            13194: color = 12'h000;
            13195: color = 12'h000;
            13196: color = 12'h000;
            13197: color = 12'h000;
            13198: color = 12'h000;
            13199: color = 12'h000;
            13200: color = 12'h000;
            13201: color = 12'h000;
            13202: color = 12'h000;
            13203: color = 12'h000;
            13204: color = 12'h000;
            13205: color = 12'h000;
            13206: color = 12'h000;
            13207: color = 12'h000;
            13208: color = 12'h000;
            13209: color = 12'h000;
            13210: color = 12'h000;
            13211: color = 12'h000;
            13212: color = 12'h000;
            13213: color = 12'h000;
            13214: color = 12'h000;
            13215: color = 12'h000;
            13216: color = 12'h000;
            13217: color = 12'h000;
            13218: color = 12'h000;
            13219: color = 12'h000;
            13220: color = 12'h000;
            13221: color = 12'h000;
            13222: color = 12'h000;
            13223: color = 12'h000;
            13224: color = 12'h000;
            13225: color = 12'h000;
            13226: color = 12'h000;
            13227: color = 12'h000;
            13228: color = 12'h000;
            13229: color = 12'h000;
            13230: color = 12'h000;
            13231: color = 12'h000;
            13232: color = 12'h000;
            13233: color = 12'h000;
            13234: color = 12'h000;
            13235: color = 12'h000;
            13236: color = 12'h000;
            13237: color = 12'h000;
            13238: color = 12'h000;
            13239: color = 12'h000;
            13240: color = 12'h000;
            13241: color = 12'h000;
            13242: color = 12'h000;
            13243: color = 12'h000;
            13244: color = 12'h000;
            13245: color = 12'h000;
            13246: color = 12'h000;
            13247: color = 12'h000;
            13248: color = 12'h000;
            13249: color = 12'h000;
            13250: color = 12'h000;
            13251: color = 12'h000;
            13252: color = 12'h000;
            13253: color = 12'h000;
            13254: color = 12'h000;
            13255: color = 12'h000;
            13256: color = 12'h000;
            13257: color = 12'h000;
            13258: color = 12'h000;
            13259: color = 12'h000;
            13260: color = 12'h000;
            13261: color = 12'h000;
            13262: color = 12'h000;
            13263: color = 12'h000;
            13264: color = 12'h000;
            13265: color = 12'h000;
            13266: color = 12'h000;
            13267: color = 12'h000;
            13268: color = 12'h000;
            13269: color = 12'h000;
            13270: color = 12'h000;
            13271: color = 12'h000;
            13272: color = 12'h000;
            13273: color = 12'h000;
            13274: color = 12'h000;
            13275: color = 12'h000;
            13276: color = 12'h000;
            13277: color = 12'h000;
            13278: color = 12'h000;
            13279: color = 12'h000;
            13280: color = 12'h000;
            13281: color = 12'h000;
            13282: color = 12'h000;
            13283: color = 12'h000;
            13284: color = 12'h000;
            13285: color = 12'h000;
            13286: color = 12'h000;
            13287: color = 12'h000;
            13288: color = 12'h000;
            13289: color = 12'h000;
            13290: color = 12'h000;
            13291: color = 12'h000;
            13292: color = 12'h000;
            13293: color = 12'h000;
            13294: color = 12'h000;
            13295: color = 12'h000;
            13296: color = 12'h000;
            13297: color = 12'h000;
            13298: color = 12'h000;
            13299: color = 12'h000;
            13300: color = 12'h000;
            13301: color = 12'h000;
            13302: color = 12'h000;
            13303: color = 12'h000;
            13304: color = 12'h000;
            13305: color = 12'h000;
            13306: color = 12'h000;
            13307: color = 12'h000;
            13308: color = 12'h000;
            13309: color = 12'h000;
            13310: color = 12'h000;
            13311: color = 12'h000;
            13312: color = 12'h000;
            13313: color = 12'h000;
            13314: color = 12'h000;
            13315: color = 12'h000;
            13316: color = 12'h000;
            13317: color = 12'h000;
            13318: color = 12'h000;
            13319: color = 12'h000;
            13320: color = 12'h000;
            13321: color = 12'h000;
            13322: color = 12'h000;
            13323: color = 12'h000;
            13324: color = 12'h000;
            13325: color = 12'h000;
            13326: color = 12'h000;
            13327: color = 12'h000;
            13328: color = 12'h000;
            13329: color = 12'h000;
            13330: color = 12'h000;
            13331: color = 12'h000;
            13332: color = 12'h000;
            13333: color = 12'h000;
            13334: color = 12'h000;
            13335: color = 12'h000;
            13336: color = 12'h000;
            13337: color = 12'h000;
            13338: color = 12'h000;
            13339: color = 12'h000;
            13340: color = 12'h000;
            13341: color = 12'h000;
            13342: color = 12'h000;
            13343: color = 12'h000;
            13344: color = 12'h000;
            13345: color = 12'h000;
            13346: color = 12'h000;
            13347: color = 12'h000;
            13348: color = 12'h000;
            13349: color = 12'h000;
            13350: color = 12'h000;
            13351: color = 12'h000;
            13352: color = 12'h000;
            13353: color = 12'h000;
            13354: color = 12'h000;
            13355: color = 12'h000;
            13356: color = 12'h000;
            13357: color = 12'h000;
            13358: color = 12'h000;
            13359: color = 12'h000;
            13360: color = 12'h000;
            13361: color = 12'h000;
            13362: color = 12'h000;
            13363: color = 12'h000;
            13364: color = 12'h000;
            13365: color = 12'h000;
            13366: color = 12'h000;
            13367: color = 12'h000;
            13368: color = 12'h000;
            13369: color = 12'h000;
            13370: color = 12'h000;
            13371: color = 12'h000;
            13372: color = 12'h000;
            13373: color = 12'h000;
            13374: color = 12'h000;
            13375: color = 12'h000;
            13376: color = 12'h000;
            13377: color = 12'h000;
            13378: color = 12'h000;
            13379: color = 12'h000;
            13380: color = 12'h000;
            13381: color = 12'h000;
            13382: color = 12'h000;
            13383: color = 12'h000;
            13384: color = 12'h000;
            13385: color = 12'h000;
            13386: color = 12'h000;
            13387: color = 12'h000;
            13388: color = 12'h000;
            13389: color = 12'h000;
            13390: color = 12'h000;
            13391: color = 12'h000;
            13392: color = 12'h000;
            13393: color = 12'h000;
            13394: color = 12'h000;
            13395: color = 12'h000;
            13396: color = 12'h000;
            13397: color = 12'h000;
            13398: color = 12'h000;
            13399: color = 12'h000;
            13400: color = 12'h000;
            13401: color = 12'h000;
            13402: color = 12'h000;
            13403: color = 12'h000;
            13404: color = 12'h000;
            13405: color = 12'h000;
            13406: color = 12'h000;
            13407: color = 12'h000;
            13408: color = 12'h000;
            13409: color = 12'h000;
            13410: color = 12'h000;
            13411: color = 12'h000;
            13412: color = 12'h000;
            13413: color = 12'h000;
            13414: color = 12'h000;
            13415: color = 12'h000;
            13416: color = 12'h000;
            13417: color = 12'h000;
            13418: color = 12'h000;
            13419: color = 12'h000;
            13420: color = 12'h000;
            13421: color = 12'h000;
            13422: color = 12'h000;
            13423: color = 12'h000;
            13424: color = 12'h000;
            13425: color = 12'h000;
            13426: color = 12'h000;
            13427: color = 12'h000;
            13428: color = 12'h000;
            13429: color = 12'h000;
            13430: color = 12'h000;
            13431: color = 12'h000;
            13432: color = 12'h000;
            13433: color = 12'h000;
            13434: color = 12'h000;
            13435: color = 12'h000;
            13436: color = 12'h000;
            13437: color = 12'h000;
            13438: color = 12'h000;
            13439: color = 12'h000;
            13440: color = 12'h000;
            13441: color = 12'h000;
            13442: color = 12'h000;
            13443: color = 12'h000;
            13444: color = 12'h000;
            13445: color = 12'h000;
            13446: color = 12'h000;
            13447: color = 12'h000;
            13448: color = 12'h000;
            13449: color = 12'h000;
            13450: color = 12'h000;
            13451: color = 12'h000;
            13452: color = 12'h000;
            13453: color = 12'h000;
            13454: color = 12'h000;
            13455: color = 12'h000;
            13456: color = 12'h000;
            13457: color = 12'h000;
            13458: color = 12'h000;
            13459: color = 12'h000;
            13460: color = 12'h000;
            13461: color = 12'h000;
            13462: color = 12'h000;
            13463: color = 12'h000;
            13464: color = 12'h000;
            13465: color = 12'h000;
            13466: color = 12'h000;
            13467: color = 12'h000;
            13468: color = 12'h000;
            13469: color = 12'h000;
            13470: color = 12'h000;
            13471: color = 12'h000;
            13472: color = 12'h000;
            13473: color = 12'h000;
            13474: color = 12'h000;
            13475: color = 12'h000;
            13476: color = 12'h000;
            13477: color = 12'h000;
            13478: color = 12'h000;
            13479: color = 12'h000;
            13480: color = 12'h000;
            13481: color = 12'h000;
            13482: color = 12'h000;
            13483: color = 12'h000;
            13484: color = 12'h000;
            13485: color = 12'h000;
            13486: color = 12'h000;
            13487: color = 12'h000;
            13488: color = 12'h000;
            13489: color = 12'h000;
            13490: color = 12'h000;
            13491: color = 12'h000;
            13492: color = 12'h000;
            13493: color = 12'h000;
            13494: color = 12'h000;
            13495: color = 12'h000;
            13496: color = 12'h000;
            13497: color = 12'h000;
            13498: color = 12'h000;
            13499: color = 12'h000;
            13500: color = 12'h000;
            13501: color = 12'h000;
            13502: color = 12'h000;
            13503: color = 12'h000;
            13504: color = 12'h000;
            13505: color = 12'h000;
            13506: color = 12'h000;
            13507: color = 12'h000;
            13508: color = 12'h000;
            13509: color = 12'h000;
            13510: color = 12'h000;
            13511: color = 12'h000;
            13512: color = 12'h000;
            13513: color = 12'h000;
            13514: color = 12'h000;
            13515: color = 12'h000;
            13516: color = 12'h000;
            13517: color = 12'h000;
            13518: color = 12'h000;
            13519: color = 12'h000;
            13520: color = 12'h000;
            13521: color = 12'h000;
            13522: color = 12'h000;
            13523: color = 12'h000;
            13524: color = 12'h000;
            13525: color = 12'h000;
            13526: color = 12'h000;
            13527: color = 12'h000;
            13528: color = 12'h000;
            13529: color = 12'h000;
            13530: color = 12'h000;
            13531: color = 12'h000;
            13532: color = 12'h000;
            13533: color = 12'h000;
            13534: color = 12'h000;
            13535: color = 12'h000;
            13536: color = 12'h000;
            13537: color = 12'h000;
            13538: color = 12'h000;
            13539: color = 12'h000;
            13540: color = 12'h000;
            13541: color = 12'h000;
            13542: color = 12'h000;
            13543: color = 12'h000;
            13544: color = 12'h000;
            13545: color = 12'h000;
            13546: color = 12'h000;
            13547: color = 12'h000;
            13548: color = 12'h000;
            13549: color = 12'h000;
            13550: color = 12'h000;
            13551: color = 12'h000;
            13552: color = 12'h000;
            13553: color = 12'h000;
            13554: color = 12'h000;
            13555: color = 12'h000;
            13556: color = 12'h000;
            13557: color = 12'h000;
            13558: color = 12'h000;
            13559: color = 12'h000;
            13560: color = 12'h000;
            13561: color = 12'h000;
            13562: color = 12'h000;
            13563: color = 12'h000;
            13564: color = 12'h000;
            13565: color = 12'h000;
            13566: color = 12'h000;
            13567: color = 12'h000;
            13568: color = 12'h000;
            13569: color = 12'h000;
            13570: color = 12'h000;
            13571: color = 12'h000;
            13572: color = 12'h000;
            13573: color = 12'h000;
            13574: color = 12'h000;
            13575: color = 12'h000;
            13576: color = 12'h000;
            13577: color = 12'h000;
            13578: color = 12'h000;
            13579: color = 12'h000;
            13580: color = 12'h000;
            13581: color = 12'h000;
            13582: color = 12'h000;
            13583: color = 12'h000;
            13584: color = 12'h000;
            13585: color = 12'h000;
            13586: color = 12'h000;
            13587: color = 12'h000;
            13588: color = 12'h000;
            13589: color = 12'h000;
            13590: color = 12'h000;
            13591: color = 12'h000;
            13592: color = 12'h000;
            13593: color = 12'h000;
            13594: color = 12'h000;
            13595: color = 12'h000;
            13596: color = 12'h000;
            13597: color = 12'h000;
            13598: color = 12'h000;
            13599: color = 12'h000;
            13600: color = 12'h000;
            13601: color = 12'h000;
            13602: color = 12'h000;
            13603: color = 12'h000;
            13604: color = 12'h000;
            13605: color = 12'h000;
            13606: color = 12'h000;
            13607: color = 12'h000;
            13608: color = 12'h000;
            13609: color = 12'h000;
            13610: color = 12'h000;
            13611: color = 12'h000;
            13612: color = 12'h000;
            13613: color = 12'h000;
            13614: color = 12'h000;
            13615: color = 12'h000;
            13616: color = 12'h000;
            13617: color = 12'h000;
            13618: color = 12'h000;
            13619: color = 12'h000;
            13620: color = 12'h000;
            13621: color = 12'h000;
            13622: color = 12'h000;
            13623: color = 12'h000;
            13624: color = 12'h000;
            13625: color = 12'h000;
            13626: color = 12'h000;
            13627: color = 12'h000;
            13628: color = 12'h000;
            13629: color = 12'h000;
            13630: color = 12'h000;
            13631: color = 12'h000;
            13632: color = 12'h000;
            13633: color = 12'h000;
            13634: color = 12'h000;
            13635: color = 12'h000;
            13636: color = 12'h000;
            13637: color = 12'h000;
            13638: color = 12'h000;
            13639: color = 12'h000;
            13640: color = 12'h000;
            13641: color = 12'h000;
            13642: color = 12'h000;
            13643: color = 12'h000;
            13644: color = 12'h000;
            13645: color = 12'h000;
            13646: color = 12'h000;
            13647: color = 12'h000;
            13648: color = 12'h000;
            13649: color = 12'h000;
            13650: color = 12'h000;
            13651: color = 12'h000;
            13652: color = 12'h000;
            13653: color = 12'h000;
            13654: color = 12'h000;
            13655: color = 12'h000;
            13656: color = 12'h000;
            13657: color = 12'h000;
            13658: color = 12'h000;
            13659: color = 12'h000;
            13660: color = 12'h000;
            13661: color = 12'h000;
            13662: color = 12'h000;
            13663: color = 12'h000;
            13664: color = 12'h000;
            13665: color = 12'h000;
            13666: color = 12'h000;
            13667: color = 12'h000;
            13668: color = 12'h000;
            13669: color = 12'h000;
            13670: color = 12'h000;
            13671: color = 12'h000;
            13672: color = 12'h000;
            13673: color = 12'h000;
            13674: color = 12'h000;
            13675: color = 12'h000;
            13676: color = 12'h000;
            13677: color = 12'h000;
            13678: color = 12'h000;
            13679: color = 12'h000;
            13680: color = 12'h000;
            13681: color = 12'h000;
            13682: color = 12'h000;
            13683: color = 12'h000;
            13684: color = 12'h000;
            13685: color = 12'h000;
            13686: color = 12'h000;
            13687: color = 12'h000;
            13688: color = 12'h000;
            13689: color = 12'h000;
            13690: color = 12'h000;
            13691: color = 12'h000;
            13692: color = 12'h000;
            13693: color = 12'h000;
            13694: color = 12'h000;
            13695: color = 12'h000;
            13696: color = 12'h000;
            13697: color = 12'h000;
            13698: color = 12'h000;
            13699: color = 12'h000;
            13700: color = 12'h000;
            13701: color = 12'h000;
            13702: color = 12'h000;
            13703: color = 12'h000;
            13704: color = 12'h000;
            13705: color = 12'h000;
            13706: color = 12'h000;
            13707: color = 12'h000;
            13708: color = 12'h000;
            13709: color = 12'h000;
            13710: color = 12'h000;
            13711: color = 12'h000;
            13712: color = 12'h000;
            13713: color = 12'h000;
            13714: color = 12'h000;
            13715: color = 12'h000;
            13716: color = 12'h000;
            13717: color = 12'h000;
            13718: color = 12'h000;
            13719: color = 12'h000;
            13720: color = 12'h000;
            13721: color = 12'h000;
            13722: color = 12'h000;
            13723: color = 12'h000;
            13724: color = 12'h000;
            13725: color = 12'h000;
            13726: color = 12'h000;
            13727: color = 12'h000;
            13728: color = 12'h000;
            13729: color = 12'h000;
            13730: color = 12'h000;
            13731: color = 12'h000;
            13732: color = 12'h000;
            13733: color = 12'h000;
            13734: color = 12'h000;
            13735: color = 12'h000;
            13736: color = 12'h000;
            13737: color = 12'h000;
            13738: color = 12'h000;
            13739: color = 12'h000;
            13740: color = 12'h000;
            13741: color = 12'h000;
            13742: color = 12'h000;
            13743: color = 12'h000;
            13744: color = 12'h000;
            13745: color = 12'h000;
            13746: color = 12'h000;
            13747: color = 12'h000;
            13748: color = 12'h000;
            13749: color = 12'h000;
            13750: color = 12'h000;
            13751: color = 12'h000;
            13752: color = 12'h000;
            13753: color = 12'h000;
            13754: color = 12'h000;
            13755: color = 12'h000;
            13756: color = 12'h000;
            13757: color = 12'h000;
            13758: color = 12'h000;
            13759: color = 12'h000;
            13760: color = 12'h000;
            13761: color = 12'h000;
            13762: color = 12'h000;
            13763: color = 12'h000;
            13764: color = 12'h000;
            13765: color = 12'h000;
            13766: color = 12'h000;
            13767: color = 12'h000;
            13768: color = 12'h000;
            13769: color = 12'h000;
            13770: color = 12'h000;
            13771: color = 12'h000;
            13772: color = 12'h000;
            13773: color = 12'h000;
            13774: color = 12'h000;
            13775: color = 12'h000;
            13776: color = 12'h000;
            13777: color = 12'h000;
            13778: color = 12'h000;
            13779: color = 12'h000;
            13780: color = 12'h000;
            13781: color = 12'h000;
            13782: color = 12'h000;
            13783: color = 12'h000;
            13784: color = 12'h000;
            13785: color = 12'h000;
            13786: color = 12'h000;
            13787: color = 12'h000;
            13788: color = 12'h000;
            13789: color = 12'h000;
            13790: color = 12'h000;
            13791: color = 12'h000;
            13792: color = 12'h000;
            13793: color = 12'h000;
            13794: color = 12'h000;
            13795: color = 12'h000;
            13796: color = 12'h000;
            13797: color = 12'h000;
            13798: color = 12'h000;
            13799: color = 12'h000;
            13800: color = 12'h000;
            13801: color = 12'h000;
            13802: color = 12'h000;
            13803: color = 12'h000;
            13804: color = 12'h000;
            13805: color = 12'h000;
            13806: color = 12'h000;
            13807: color = 12'h000;
            13808: color = 12'h000;
            13809: color = 12'h000;
            13810: color = 12'h000;
            13811: color = 12'h000;
            13812: color = 12'h000;
            13813: color = 12'h000;
            13814: color = 12'h000;
            13815: color = 12'h000;
            13816: color = 12'h000;
            13817: color = 12'h000;
            13818: color = 12'h000;
            13819: color = 12'h000;
            13820: color = 12'h000;
            13821: color = 12'h000;
            13822: color = 12'h000;
            13823: color = 12'h000;
            13824: color = 12'h000;
            13825: color = 12'h000;
            13826: color = 12'h000;
            13827: color = 12'h000;
            13828: color = 12'h000;
            13829: color = 12'h000;
            13830: color = 12'h000;
            13831: color = 12'h000;
            13832: color = 12'h000;
            13833: color = 12'h000;
            13834: color = 12'h000;
            13835: color = 12'h000;
            13836: color = 12'h000;
            13837: color = 12'h000;
            13838: color = 12'h000;
            13839: color = 12'h000;
            13840: color = 12'h000;
            13841: color = 12'h000;
            13842: color = 12'h000;
            13843: color = 12'h000;
            13844: color = 12'h000;
            13845: color = 12'h000;
            13846: color = 12'h000;
            13847: color = 12'h000;
            13848: color = 12'h000;
            13849: color = 12'h000;
            13850: color = 12'h000;
            13851: color = 12'h000;
            13852: color = 12'h000;
            13853: color = 12'h000;
            13854: color = 12'h000;
            13855: color = 12'h000;
            13856: color = 12'h000;
            13857: color = 12'h000;
            13858: color = 12'h000;
            13859: color = 12'h000;
            13860: color = 12'h000;
            13861: color = 12'h000;
            13862: color = 12'h000;
            13863: color = 12'h000;
            13864: color = 12'h000;
            13865: color = 12'h000;
            13866: color = 12'h000;
            13867: color = 12'h000;
            13868: color = 12'h000;
            13869: color = 12'h000;
            13870: color = 12'h000;
            13871: color = 12'h000;
            13872: color = 12'h000;
            13873: color = 12'h000;
            13874: color = 12'h000;
            13875: color = 12'h000;
            13876: color = 12'h000;
            13877: color = 12'h000;
            13878: color = 12'h000;
            13879: color = 12'h000;
            13880: color = 12'h000;
            13881: color = 12'h000;
            13882: color = 12'h000;
            13883: color = 12'h000;
            13884: color = 12'h000;
            13885: color = 12'h000;
            13886: color = 12'h000;
            13887: color = 12'h000;
            13888: color = 12'h000;
            13889: color = 12'h000;
            13890: color = 12'h000;
            13891: color = 12'h000;
            13892: color = 12'h000;
            13893: color = 12'h000;
            13894: color = 12'h000;
            13895: color = 12'h000;
            13896: color = 12'h000;
            13897: color = 12'h000;
            13898: color = 12'h000;
            13899: color = 12'h000;
            13900: color = 12'h000;
            13901: color = 12'h000;
            13902: color = 12'h000;
            13903: color = 12'h000;
            13904: color = 12'h000;
            13905: color = 12'h000;
            13906: color = 12'h000;
            13907: color = 12'h000;
            13908: color = 12'h000;
            13909: color = 12'h000;
            13910: color = 12'h000;
            13911: color = 12'h000;
            13912: color = 12'h000;
            13913: color = 12'h000;
            13914: color = 12'h000;
            13915: color = 12'h000;
            13916: color = 12'h000;
            13917: color = 12'h000;
            13918: color = 12'h000;
            13919: color = 12'h000;
            13920: color = 12'h000;
            13921: color = 12'h000;
            13922: color = 12'h000;
            13923: color = 12'h000;
            13924: color = 12'h000;
            13925: color = 12'h000;
            13926: color = 12'h000;
            13927: color = 12'h000;
            13928: color = 12'h000;
            13929: color = 12'h000;
            13930: color = 12'h000;
            13931: color = 12'h000;
            13932: color = 12'h000;
            13933: color = 12'h000;
            13934: color = 12'h000;
            13935: color = 12'h000;
            13936: color = 12'h000;
            13937: color = 12'h000;
            13938: color = 12'h000;
            13939: color = 12'h000;
            13940: color = 12'h000;
            13941: color = 12'h000;
            13942: color = 12'h000;
            13943: color = 12'h000;
            13944: color = 12'h000;
            13945: color = 12'h000;
            13946: color = 12'h000;
            13947: color = 12'h000;
            13948: color = 12'h000;
            13949: color = 12'h000;
            13950: color = 12'h000;
            13951: color = 12'h000;
            13952: color = 12'h000;
            13953: color = 12'h000;
            13954: color = 12'h000;
            13955: color = 12'h000;
            13956: color = 12'h000;
            13957: color = 12'h000;
            13958: color = 12'h000;
            13959: color = 12'h000;
            13960: color = 12'h000;
            13961: color = 12'h000;
            13962: color = 12'h000;
            13963: color = 12'h000;
            13964: color = 12'h000;
            13965: color = 12'h000;
            13966: color = 12'h000;
            13967: color = 12'h000;
            13968: color = 12'h000;
            13969: color = 12'h000;
            13970: color = 12'h000;
            13971: color = 12'h000;
            13972: color = 12'h000;
            13973: color = 12'h000;
            13974: color = 12'h000;
            13975: color = 12'h000;
            13976: color = 12'h000;
            13977: color = 12'h000;
            13978: color = 12'h000;
            13979: color = 12'h000;
            13980: color = 12'h000;
            13981: color = 12'h000;
            13982: color = 12'h000;
            13983: color = 12'h000;
            13984: color = 12'h000;
            13985: color = 12'h000;
            13986: color = 12'h000;
            13987: color = 12'h000;
            13988: color = 12'h000;
            13989: color = 12'h000;
            13990: color = 12'h000;
            13991: color = 12'h000;
            13992: color = 12'h000;
            13993: color = 12'h000;
            13994: color = 12'h000;
            13995: color = 12'h000;
            13996: color = 12'h000;
            13997: color = 12'h000;
            13998: color = 12'h000;
            13999: color = 12'h000;
            14000: color = 12'h000;
            14001: color = 12'h000;
            14002: color = 12'h000;
            14003: color = 12'h000;
            14004: color = 12'h000;
            14005: color = 12'h000;
            14006: color = 12'h000;
            14007: color = 12'h000;
            14008: color = 12'h000;
            14009: color = 12'h000;
            14010: color = 12'h000;
            14011: color = 12'h000;
            14012: color = 12'h000;
            14013: color = 12'h000;
            14014: color = 12'h000;
            14015: color = 12'h000;
            14016: color = 12'h000;
            14017: color = 12'h000;
            14018: color = 12'h000;
            14019: color = 12'h000;
            14020: color = 12'h000;
            14021: color = 12'h000;
            14022: color = 12'h000;
            14023: color = 12'h000;
            14024: color = 12'h000;
            14025: color = 12'h000;
            14026: color = 12'h000;
            14027: color = 12'h000;
            14028: color = 12'h000;
            14029: color = 12'h000;
            14030: color = 12'h000;
            14031: color = 12'h000;
            14032: color = 12'h000;
            14033: color = 12'h000;
            14034: color = 12'h000;
            14035: color = 12'h000;
            14036: color = 12'h000;
            14037: color = 12'h000;
            14038: color = 12'h000;
            14039: color = 12'h000;
            14040: color = 12'h000;
            14041: color = 12'h000;
            14042: color = 12'h000;
            14043: color = 12'h000;
            14044: color = 12'h000;
            14045: color = 12'h000;
            14046: color = 12'h000;
            14047: color = 12'h000;
            14048: color = 12'h000;
            14049: color = 12'h000;
            14050: color = 12'h000;
            14051: color = 12'h000;
            14052: color = 12'h000;
            14053: color = 12'h000;
            14054: color = 12'h000;
            14055: color = 12'h000;
            14056: color = 12'h000;
            14057: color = 12'h000;
            14058: color = 12'h000;
            14059: color = 12'h000;
            14060: color = 12'h000;
            14061: color = 12'h000;
            14062: color = 12'h000;
            14063: color = 12'h000;
            14064: color = 12'h000;
            14065: color = 12'h000;
            14066: color = 12'h000;
            14067: color = 12'h000;
            14068: color = 12'h000;
            14069: color = 12'h000;
            14070: color = 12'h000;
            14071: color = 12'h000;
            14072: color = 12'h000;
            14073: color = 12'h000;
            14074: color = 12'h000;
            14075: color = 12'h000;
            14076: color = 12'h000;
            14077: color = 12'h000;
            14078: color = 12'h000;
            14079: color = 12'h000;
            14080: color = 12'h000;
            14081: color = 12'h000;
            14082: color = 12'h000;
            14083: color = 12'h000;
            14084: color = 12'h000;
            14085: color = 12'h000;
            14086: color = 12'h000;
            14087: color = 12'h000;
            14088: color = 12'h000;
            14089: color = 12'h000;
            14090: color = 12'h000;
            14091: color = 12'h000;
            14092: color = 12'h000;
            14093: color = 12'h000;
            14094: color = 12'h000;
            14095: color = 12'h000;
            14096: color = 12'h000;
            14097: color = 12'h000;
            14098: color = 12'h000;
            14099: color = 12'h000;
            14100: color = 12'h000;
            14101: color = 12'h000;
            14102: color = 12'h000;
            14103: color = 12'h000;
            14104: color = 12'h000;
            14105: color = 12'h000;
            14106: color = 12'h000;
            14107: color = 12'h000;
            14108: color = 12'h000;
            14109: color = 12'h000;
            14110: color = 12'h000;
            14111: color = 12'h000;
            14112: color = 12'h000;
            14113: color = 12'h000;
            14114: color = 12'h000;
            14115: color = 12'h000;
            14116: color = 12'h000;
            14117: color = 12'h000;
            14118: color = 12'h000;
            14119: color = 12'h000;
            14120: color = 12'h000;
            14121: color = 12'h000;
            14122: color = 12'h000;
            14123: color = 12'h000;
            14124: color = 12'h000;
            14125: color = 12'h000;
            14126: color = 12'h000;
            14127: color = 12'h000;
            14128: color = 12'h000;
            14129: color = 12'h000;
            14130: color = 12'h000;
            14131: color = 12'h000;
            14132: color = 12'h000;
            14133: color = 12'h000;
            14134: color = 12'h000;
            14135: color = 12'h000;
            14136: color = 12'h000;
            14137: color = 12'h000;
            14138: color = 12'h000;
            14139: color = 12'h000;
            14140: color = 12'h000;
            14141: color = 12'h000;
            14142: color = 12'h000;
            14143: color = 12'h000;
            14144: color = 12'h000;
            14145: color = 12'h000;
            14146: color = 12'h000;
            14147: color = 12'h000;
            14148: color = 12'h000;
            14149: color = 12'h000;
            14150: color = 12'h000;
            14151: color = 12'h000;
            14152: color = 12'h000;
            14153: color = 12'h000;
            14154: color = 12'h000;
            14155: color = 12'h000;
            14156: color = 12'h000;
            14157: color = 12'h000;
            14158: color = 12'h000;
            14159: color = 12'h000;
            14160: color = 12'h000;
            14161: color = 12'h000;
            14162: color = 12'h000;
            14163: color = 12'h000;
            14164: color = 12'h000;
            14165: color = 12'h000;
            14166: color = 12'h000;
            14167: color = 12'h000;
            14168: color = 12'h000;
            14169: color = 12'h000;
            14170: color = 12'h000;
            14171: color = 12'h000;
            14172: color = 12'h000;
            14173: color = 12'h000;
            14174: color = 12'h000;
            14175: color = 12'h000;
            14176: color = 12'h000;
            14177: color = 12'h000;
            14178: color = 12'h000;
            14179: color = 12'h000;
            14180: color = 12'h000;
            14181: color = 12'h000;
            14182: color = 12'h000;
            14183: color = 12'h000;
            14184: color = 12'h000;
            14185: color = 12'h000;
            14186: color = 12'h000;
            14187: color = 12'h000;
            14188: color = 12'h000;
            14189: color = 12'h000;
            14190: color = 12'h000;
            14191: color = 12'h000;
            14192: color = 12'h000;
            14193: color = 12'h000;
            14194: color = 12'h000;
            14195: color = 12'h000;
            14196: color = 12'h000;
            14197: color = 12'h000;
            14198: color = 12'h000;
            14199: color = 12'h000;
            14200: color = 12'h000;
            14201: color = 12'h000;
            14202: color = 12'h000;
            14203: color = 12'h000;
            14204: color = 12'h000;
            14205: color = 12'h000;
            14206: color = 12'h000;
            14207: color = 12'h000;
            14208: color = 12'h000;
            14209: color = 12'h000;
            14210: color = 12'h000;
            14211: color = 12'h000;
            14212: color = 12'h000;
            14213: color = 12'h000;
            14214: color = 12'h000;
            14215: color = 12'h000;
            14216: color = 12'h000;
            14217: color = 12'h000;
            14218: color = 12'h000;
            14219: color = 12'h000;
            14220: color = 12'h000;
            14221: color = 12'h000;
            14222: color = 12'h000;
            14223: color = 12'h000;
            14224: color = 12'h000;
            14225: color = 12'h000;
            14226: color = 12'h000;
            14227: color = 12'h000;
            14228: color = 12'h000;
            14229: color = 12'h000;
            14230: color = 12'h000;
            14231: color = 12'h000;
            14232: color = 12'h000;
            14233: color = 12'h000;
            14234: color = 12'h000;
            14235: color = 12'h000;
            14236: color = 12'h000;
            14237: color = 12'h000;
            14238: color = 12'h000;
            14239: color = 12'h000;
            14240: color = 12'h000;
            14241: color = 12'h000;
            14242: color = 12'h000;
            14243: color = 12'h000;
            14244: color = 12'h000;
            14245: color = 12'h000;
            14246: color = 12'h000;
            14247: color = 12'h000;
            14248: color = 12'h000;
            14249: color = 12'h000;
            14250: color = 12'h000;
            14251: color = 12'h000;
            14252: color = 12'h000;
            14253: color = 12'h000;
            14254: color = 12'h000;
            14255: color = 12'h000;
            14256: color = 12'h000;
            14257: color = 12'h000;
            14258: color = 12'h000;
            14259: color = 12'h000;
            14260: color = 12'h000;
            14261: color = 12'h000;
            14262: color = 12'h000;
            14263: color = 12'h000;
            14264: color = 12'h000;
            14265: color = 12'h000;
            14266: color = 12'h000;
            14267: color = 12'h000;
            14268: color = 12'h000;
            14269: color = 12'h000;
            14270: color = 12'h000;
            14271: color = 12'h000;
            14272: color = 12'h000;
            14273: color = 12'h000;
            14274: color = 12'h000;
            14275: color = 12'h000;
            14276: color = 12'h000;
            14277: color = 12'h000;
            14278: color = 12'h000;
            14279: color = 12'h000;
            14280: color = 12'h000;
            14281: color = 12'h000;
            14282: color = 12'h000;
            14283: color = 12'h000;
            14284: color = 12'h000;
            14285: color = 12'h000;
            14286: color = 12'h000;
            14287: color = 12'h000;
            14288: color = 12'h000;
            14289: color = 12'h000;
            14290: color = 12'h000;
            14291: color = 12'h000;
            14292: color = 12'h000;
            14293: color = 12'h000;
            14294: color = 12'h000;
            14295: color = 12'h000;
            14296: color = 12'h000;
            14297: color = 12'h000;
            14298: color = 12'h000;
            14299: color = 12'h000;
            14300: color = 12'h000;
            14301: color = 12'h000;
            14302: color = 12'h000;
            14303: color = 12'h000;
            14304: color = 12'h000;
            14305: color = 12'h000;
            14306: color = 12'h000;
            14307: color = 12'h000;
            14308: color = 12'h000;
            14309: color = 12'h000;
            14310: color = 12'h000;
            14311: color = 12'h000;
            14312: color = 12'h000;
            14313: color = 12'h000;
            14314: color = 12'h000;
            14315: color = 12'h000;
            14316: color = 12'h000;
            14317: color = 12'h000;
            14318: color = 12'h000;
            14319: color = 12'h000;
            14320: color = 12'h000;
            14321: color = 12'h000;
            14322: color = 12'h000;
            14323: color = 12'h000;
            14324: color = 12'h000;
            14325: color = 12'h000;
            14326: color = 12'h000;
            14327: color = 12'h000;
            14328: color = 12'h000;
            14329: color = 12'h000;
            14330: color = 12'h000;
            14331: color = 12'h000;
            14332: color = 12'h000;
            14333: color = 12'h000;
            14334: color = 12'h000;
            14335: color = 12'h000;
            14336: color = 12'h000;
            14337: color = 12'h000;
            14338: color = 12'h000;
            14339: color = 12'h000;
            14340: color = 12'h000;
            14341: color = 12'h000;
            14342: color = 12'h000;
            14343: color = 12'h000;
            14344: color = 12'h000;
            14345: color = 12'h000;
            14346: color = 12'h000;
            14347: color = 12'h000;
            14348: color = 12'h000;
            14349: color = 12'h000;
            14350: color = 12'h000;
            14351: color = 12'h000;
            14352: color = 12'h000;
            14353: color = 12'h000;
            14354: color = 12'h000;
            14355: color = 12'h000;
            14356: color = 12'h000;
            14357: color = 12'h000;
            14358: color = 12'h000;
            14359: color = 12'h000;
            14360: color = 12'h000;
            14361: color = 12'h000;
            14362: color = 12'h000;
            14363: color = 12'h000;
            14364: color = 12'h000;
            14365: color = 12'h000;
            14366: color = 12'h000;
            14367: color = 12'h000;
            14368: color = 12'h000;
            14369: color = 12'h000;
            14370: color = 12'h000;
            14371: color = 12'h000;
            14372: color = 12'h000;
            14373: color = 12'h000;
            14374: color = 12'h000;
            14375: color = 12'h000;
            14376: color = 12'h000;
            14377: color = 12'h000;
            14378: color = 12'h000;
            14379: color = 12'h000;
            14380: color = 12'h000;
            14381: color = 12'h000;
            14382: color = 12'h000;
            14383: color = 12'h000;
            14384: color = 12'h000;
            14385: color = 12'h000;
            14386: color = 12'h000;
            14387: color = 12'h000;
            14388: color = 12'h000;
            14389: color = 12'h000;
            14390: color = 12'h000;
            14391: color = 12'h000;
            14392: color = 12'h000;
            14393: color = 12'h000;
            14394: color = 12'h000;
            14395: color = 12'h000;
            14396: color = 12'h000;
            14397: color = 12'h000;
            14398: color = 12'h000;
            14399: color = 12'h000;
            14400: color = 12'h000;
            14401: color = 12'h000;
            14402: color = 12'h000;
            14403: color = 12'h000;
            14404: color = 12'h000;
            14405: color = 12'h000;
            14406: color = 12'h000;
            14407: color = 12'h000;
            14408: color = 12'h000;
            14409: color = 12'h000;
            14410: color = 12'h000;
            14411: color = 12'h000;
            14412: color = 12'h000;
            14413: color = 12'h000;
            14414: color = 12'h000;
            14415: color = 12'h000;
            14416: color = 12'h000;
            14417: color = 12'h000;
            14418: color = 12'h000;
            14419: color = 12'h000;
            14420: color = 12'h000;
            14421: color = 12'h000;
            14422: color = 12'h000;
            14423: color = 12'h000;
            14424: color = 12'h000;
            14425: color = 12'h000;
            14426: color = 12'h000;
            14427: color = 12'h000;
            14428: color = 12'h000;
            14429: color = 12'h000;
            14430: color = 12'h000;
            14431: color = 12'h000;
            14432: color = 12'h000;
            14433: color = 12'h000;
            14434: color = 12'h000;
            14435: color = 12'h000;
            14436: color = 12'h000;
            14437: color = 12'h000;
            14438: color = 12'h000;
            14439: color = 12'h000;
            14440: color = 12'h000;
            14441: color = 12'h000;
            14442: color = 12'h000;
            14443: color = 12'h000;
            14444: color = 12'h000;
            14445: color = 12'h000;
            14446: color = 12'h000;
            14447: color = 12'h000;
            14448: color = 12'h000;
            14449: color = 12'h000;
            14450: color = 12'h000;
            14451: color = 12'h000;
            14452: color = 12'h000;
            14453: color = 12'h000;
            14454: color = 12'h000;
            14455: color = 12'h000;
            14456: color = 12'h000;
            14457: color = 12'h000;
            14458: color = 12'h000;
            14459: color = 12'h000;
            14460: color = 12'h000;
            14461: color = 12'h000;
            14462: color = 12'h000;
            14463: color = 12'h000;
            14464: color = 12'h000;
            14465: color = 12'h000;
            14466: color = 12'h000;
            14467: color = 12'h000;
            14468: color = 12'h000;
            14469: color = 12'h000;
            14470: color = 12'h000;
            14471: color = 12'h000;
            14472: color = 12'h000;
            14473: color = 12'h000;
            14474: color = 12'h000;
            14475: color = 12'h000;
            14476: color = 12'h000;
            14477: color = 12'h000;
            14478: color = 12'h000;
            14479: color = 12'h000;
            14480: color = 12'h000;
            14481: color = 12'h000;
            14482: color = 12'h000;
            14483: color = 12'h000;
            14484: color = 12'h000;
            14485: color = 12'h000;
            14486: color = 12'h000;
            14487: color = 12'h000;
            14488: color = 12'h000;
            14489: color = 12'h000;
            14490: color = 12'h000;
            14491: color = 12'h000;
            14492: color = 12'h000;
            14493: color = 12'h000;
            14494: color = 12'h000;
            14495: color = 12'h000;
            14496: color = 12'h000;
            14497: color = 12'h000;
            14498: color = 12'h000;
            14499: color = 12'h000;
            14500: color = 12'h000;
            14501: color = 12'h000;
            14502: color = 12'h000;
            14503: color = 12'h000;
            14504: color = 12'h000;
            14505: color = 12'h000;
            14506: color = 12'h000;
            14507: color = 12'h000;
            14508: color = 12'h000;
            14509: color = 12'h000;
            14510: color = 12'h000;
            14511: color = 12'h000;
            14512: color = 12'h000;
            14513: color = 12'h000;
            14514: color = 12'h000;
            14515: color = 12'h000;
            14516: color = 12'h000;
            14517: color = 12'h000;
            14518: color = 12'h000;
            14519: color = 12'h000;
            14520: color = 12'h000;
            14521: color = 12'h000;
            14522: color = 12'h000;
            14523: color = 12'h000;
            14524: color = 12'h000;
            14525: color = 12'h000;
            14526: color = 12'h000;
            14527: color = 12'h000;
            14528: color = 12'h000;
            14529: color = 12'h000;
            14530: color = 12'h000;
            14531: color = 12'h000;
            14532: color = 12'h000;
            14533: color = 12'h000;
            14534: color = 12'h000;
            14535: color = 12'h000;
            14536: color = 12'h000;
            14537: color = 12'h000;
            14538: color = 12'h000;
            14539: color = 12'h000;
            14540: color = 12'h000;
            14541: color = 12'h000;
            14542: color = 12'h000;
            14543: color = 12'h000;
            14544: color = 12'h000;
            14545: color = 12'h000;
            14546: color = 12'h000;
            14547: color = 12'h000;
            14548: color = 12'h000;
            14549: color = 12'h000;
            14550: color = 12'h000;
            14551: color = 12'h000;
            14552: color = 12'h000;
            14553: color = 12'h000;
            14554: color = 12'h000;
            14555: color = 12'h000;
            14556: color = 12'h000;
            14557: color = 12'h000;
            14558: color = 12'h000;
            14559: color = 12'h000;
            14560: color = 12'h000;
            14561: color = 12'h000;
            14562: color = 12'h000;
            14563: color = 12'h000;
            14564: color = 12'h000;
            14565: color = 12'h000;
            14566: color = 12'h000;
            14567: color = 12'h000;
            14568: color = 12'h000;
            14569: color = 12'h000;
            14570: color = 12'h000;
            14571: color = 12'h000;
            14572: color = 12'h000;
            14573: color = 12'h000;
            14574: color = 12'h000;
            14575: color = 12'h000;
            14576: color = 12'h000;
            14577: color = 12'h000;
            14578: color = 12'h000;
            14579: color = 12'h000;
            14580: color = 12'h000;
            14581: color = 12'h000;
            14582: color = 12'h000;
            14583: color = 12'h000;
            14584: color = 12'h000;
            14585: color = 12'h000;
            14586: color = 12'h000;
            14587: color = 12'h000;
            14588: color = 12'h000;
            14589: color = 12'h000;
            14590: color = 12'h000;
            14591: color = 12'h000;
            14592: color = 12'h000;
            14593: color = 12'h000;
            14594: color = 12'h000;
            14595: color = 12'h000;
            14596: color = 12'h000;
            14597: color = 12'h000;
            14598: color = 12'h000;
            14599: color = 12'h000;
            14600: color = 12'h000;
            14601: color = 12'h000;
            14602: color = 12'h000;
            14603: color = 12'h000;
            14604: color = 12'h000;
            14605: color = 12'h000;
            14606: color = 12'h000;
            14607: color = 12'h000;
            14608: color = 12'h000;
            14609: color = 12'h000;
            14610: color = 12'h000;
            14611: color = 12'h000;
            14612: color = 12'h000;
            14613: color = 12'h000;
            14614: color = 12'h000;
            14615: color = 12'h000;
            14616: color = 12'h000;
            14617: color = 12'h000;
            14618: color = 12'h000;
            14619: color = 12'h000;
            14620: color = 12'h000;
            14621: color = 12'h000;
            14622: color = 12'h000;
            14623: color = 12'h000;
            14624: color = 12'h000;
            14625: color = 12'h000;
            14626: color = 12'h000;
            14627: color = 12'h000;
            14628: color = 12'h000;
            14629: color = 12'h000;
            14630: color = 12'h000;
            14631: color = 12'h000;
            14632: color = 12'h000;
            14633: color = 12'h000;
            14634: color = 12'h000;
            14635: color = 12'h000;
            14636: color = 12'h000;
            14637: color = 12'h000;
            14638: color = 12'h000;
            14639: color = 12'h000;
            14640: color = 12'h000;
            14641: color = 12'h000;
            14642: color = 12'h000;
            14643: color = 12'h000;
            14644: color = 12'h000;
            14645: color = 12'h000;
            14646: color = 12'h000;
            14647: color = 12'h000;
            14648: color = 12'h000;
            14649: color = 12'h000;
            14650: color = 12'h000;
            14651: color = 12'h000;
            14652: color = 12'h000;
            14653: color = 12'h000;
            14654: color = 12'h000;
            14655: color = 12'h000;
            14656: color = 12'h000;
            14657: color = 12'h000;
            14658: color = 12'h000;
            14659: color = 12'h000;
            14660: color = 12'h000;
            14661: color = 12'h000;
            14662: color = 12'h000;
            14663: color = 12'h000;
            14664: color = 12'h000;
            14665: color = 12'h000;
            14666: color = 12'h000;
            14667: color = 12'h000;
            14668: color = 12'h000;
            14669: color = 12'h000;
            14670: color = 12'h000;
            14671: color = 12'h000;
            14672: color = 12'h000;
            14673: color = 12'h000;
            14674: color = 12'h000;
            14675: color = 12'h000;
            14676: color = 12'h000;
            14677: color = 12'h000;
            14678: color = 12'h000;
            14679: color = 12'h000;
            14680: color = 12'h000;
            14681: color = 12'h000;
            14682: color = 12'h000;
            14683: color = 12'h000;
            14684: color = 12'h000;
            14685: color = 12'h000;
            14686: color = 12'h000;
            14687: color = 12'h000;
            14688: color = 12'h000;
            14689: color = 12'h000;
            14690: color = 12'h000;
            14691: color = 12'h000;
            14692: color = 12'h000;
            14693: color = 12'h000;
            14694: color = 12'h000;
            14695: color = 12'h000;
            14696: color = 12'h000;
            14697: color = 12'h000;
            14698: color = 12'h000;
            14699: color = 12'h000;
            14700: color = 12'h000;
            14701: color = 12'h000;
            14702: color = 12'h000;
            14703: color = 12'h000;
            14704: color = 12'h000;
            14705: color = 12'h000;
            14706: color = 12'h000;
            14707: color = 12'h000;
            14708: color = 12'h000;
            14709: color = 12'h000;
            14710: color = 12'h000;
            14711: color = 12'h000;
            14712: color = 12'h000;
            14713: color = 12'h000;
            14714: color = 12'h000;
            14715: color = 12'h000;
            14716: color = 12'h000;
            14717: color = 12'h000;
            14718: color = 12'h000;
            14719: color = 12'h000;
            14720: color = 12'h000;
            14721: color = 12'h000;
            14722: color = 12'h000;
            14723: color = 12'h000;
            14724: color = 12'h000;
            14725: color = 12'h000;
            14726: color = 12'h000;
            14727: color = 12'h000;
            14728: color = 12'h000;
            14729: color = 12'h000;
            14730: color = 12'h000;
            14731: color = 12'h000;
            14732: color = 12'h000;
            14733: color = 12'h000;
            14734: color = 12'h000;
            14735: color = 12'h000;
            14736: color = 12'h000;
            14737: color = 12'h000;
            14738: color = 12'h000;
            14739: color = 12'h000;
            14740: color = 12'h000;
            14741: color = 12'h000;
            14742: color = 12'h000;
            14743: color = 12'h000;
            14744: color = 12'h000;
            14745: color = 12'h000;
            14746: color = 12'h000;
            14747: color = 12'h000;
            14748: color = 12'h000;
            14749: color = 12'h000;
            14750: color = 12'h000;
            14751: color = 12'h000;
            14752: color = 12'h000;
            14753: color = 12'h000;
            14754: color = 12'h000;
            14755: color = 12'h000;
            14756: color = 12'h000;
            14757: color = 12'h000;
            14758: color = 12'h000;
            14759: color = 12'h000;
            14760: color = 12'h000;
            14761: color = 12'h000;
            14762: color = 12'h000;
            14763: color = 12'h000;
            14764: color = 12'h000;
            14765: color = 12'h000;
            14766: color = 12'h000;
            14767: color = 12'h000;
            14768: color = 12'h000;
            14769: color = 12'h000;
            14770: color = 12'h000;
            14771: color = 12'h000;
            14772: color = 12'h000;
            14773: color = 12'h000;
            14774: color = 12'h000;
            14775: color = 12'h000;
            14776: color = 12'h000;
            14777: color = 12'h000;
            14778: color = 12'h000;
            14779: color = 12'h000;
            14780: color = 12'h000;
            14781: color = 12'h000;
            14782: color = 12'h000;
            14783: color = 12'h000;
            14784: color = 12'h000;
            14785: color = 12'h000;
            14786: color = 12'h000;
            14787: color = 12'h000;
            14788: color = 12'h000;
            14789: color = 12'h000;
            14790: color = 12'h000;
            14791: color = 12'h000;
            14792: color = 12'h000;
            14793: color = 12'h000;
            14794: color = 12'h000;
            14795: color = 12'h000;
            14796: color = 12'h000;
            14797: color = 12'h000;
            14798: color = 12'h000;
            14799: color = 12'h000;
            14800: color = 12'h000;
            14801: color = 12'h000;
            14802: color = 12'h000;
            14803: color = 12'h000;
            14804: color = 12'h000;
            14805: color = 12'h000;
            14806: color = 12'h000;
            14807: color = 12'h000;
            14808: color = 12'h000;
            14809: color = 12'h000;
            14810: color = 12'h000;
            14811: color = 12'h000;
            14812: color = 12'h000;
            14813: color = 12'h000;
            14814: color = 12'h000;
            14815: color = 12'h000;
            14816: color = 12'h000;
            14817: color = 12'h000;
            14818: color = 12'h000;
            14819: color = 12'h000;
            14820: color = 12'h000;
            14821: color = 12'h000;
            14822: color = 12'h000;
            14823: color = 12'h000;
            14824: color = 12'h000;
            14825: color = 12'h000;
            14826: color = 12'h000;
            14827: color = 12'h000;
            14828: color = 12'h000;
            14829: color = 12'h000;
            14830: color = 12'h000;
            14831: color = 12'h000;
            14832: color = 12'h000;
            14833: color = 12'h000;
            14834: color = 12'h000;
            14835: color = 12'h000;
            14836: color = 12'h000;
            14837: color = 12'h000;
            14838: color = 12'h000;
            14839: color = 12'h000;
            14840: color = 12'h000;
            14841: color = 12'h000;
            14842: color = 12'h000;
            14843: color = 12'h000;
            14844: color = 12'h000;
            14845: color = 12'h000;
            14846: color = 12'h000;
            14847: color = 12'h000;
            14848: color = 12'h000;
            14849: color = 12'h000;
            14850: color = 12'h000;
            14851: color = 12'h000;
            14852: color = 12'h000;
            14853: color = 12'h000;
            14854: color = 12'h000;
            14855: color = 12'h000;
            14856: color = 12'h000;
            14857: color = 12'h000;
            14858: color = 12'h000;
            14859: color = 12'h000;
            14860: color = 12'h000;
            14861: color = 12'h000;
            14862: color = 12'h000;
            14863: color = 12'h000;
            14864: color = 12'h000;
            14865: color = 12'h000;
            14866: color = 12'h000;
            14867: color = 12'h000;
            14868: color = 12'h000;
            14869: color = 12'h000;
            14870: color = 12'h000;
            14871: color = 12'h000;
            14872: color = 12'h000;
            14873: color = 12'h000;
            14874: color = 12'h000;
            14875: color = 12'h000;
            14876: color = 12'h000;
            14877: color = 12'h000;
            14878: color = 12'h000;
            14879: color = 12'h000;
            14880: color = 12'h000;
            14881: color = 12'h000;
            14882: color = 12'h000;
            14883: color = 12'h000;
            14884: color = 12'h000;
            14885: color = 12'h000;
            14886: color = 12'h000;
            14887: color = 12'h000;
            14888: color = 12'h000;
            14889: color = 12'h000;
            14890: color = 12'h000;
            14891: color = 12'h000;
            14892: color = 12'h000;
            14893: color = 12'h000;
            14894: color = 12'h000;
            14895: color = 12'h000;
            14896: color = 12'h000;
            14897: color = 12'h000;
            14898: color = 12'h000;
            14899: color = 12'h000;
            14900: color = 12'h000;
            14901: color = 12'h000;
            14902: color = 12'h000;
            14903: color = 12'h000;
            14904: color = 12'h000;
            14905: color = 12'h000;
            14906: color = 12'h000;
            14907: color = 12'h000;
            14908: color = 12'h000;
            14909: color = 12'h000;
            14910: color = 12'h000;
            14911: color = 12'h000;
            14912: color = 12'h000;
            14913: color = 12'h000;
            14914: color = 12'h000;
            14915: color = 12'h000;
            14916: color = 12'h000;
            14917: color = 12'h000;
            14918: color = 12'h000;
            14919: color = 12'h000;
            14920: color = 12'h000;
            14921: color = 12'h000;
            14922: color = 12'h000;
            14923: color = 12'h000;
            14924: color = 12'h000;
            14925: color = 12'h000;
            14926: color = 12'h000;
            14927: color = 12'h000;
            14928: color = 12'h000;
            14929: color = 12'h000;
            14930: color = 12'h000;
            14931: color = 12'h000;
            14932: color = 12'h000;
            14933: color = 12'h000;
            14934: color = 12'h000;
            14935: color = 12'h000;
            14936: color = 12'h000;
            14937: color = 12'h000;
            14938: color = 12'h000;
            14939: color = 12'h000;
            14940: color = 12'h000;
            14941: color = 12'h000;
            14942: color = 12'h000;
            14943: color = 12'h000;
            14944: color = 12'h000;
            14945: color = 12'h000;
            14946: color = 12'h000;
            14947: color = 12'h000;
            14948: color = 12'h000;
            14949: color = 12'h000;
            14950: color = 12'h000;
            14951: color = 12'h000;
            14952: color = 12'h000;
            14953: color = 12'h000;
            14954: color = 12'h000;
            14955: color = 12'h000;
            14956: color = 12'h000;
            14957: color = 12'h000;
            14958: color = 12'h000;
            14959: color = 12'h000;
            14960: color = 12'h000;
            14961: color = 12'h000;
            14962: color = 12'h000;
            14963: color = 12'h000;
            14964: color = 12'h000;
            14965: color = 12'h000;
            14966: color = 12'h000;
            14967: color = 12'h000;
            14968: color = 12'h000;
            14969: color = 12'h000;
            14970: color = 12'h000;
            14971: color = 12'h000;
            14972: color = 12'h000;
            14973: color = 12'h000;
            14974: color = 12'h000;
            14975: color = 12'h000;
            14976: color = 12'h000;
            14977: color = 12'h000;
            14978: color = 12'h000;
            14979: color = 12'h000;
            14980: color = 12'h000;
            14981: color = 12'h000;
            14982: color = 12'h000;
            14983: color = 12'h000;
            14984: color = 12'h000;
            14985: color = 12'h000;
            14986: color = 12'h000;
            14987: color = 12'h000;
            14988: color = 12'h000;
            14989: color = 12'h000;
            14990: color = 12'h000;
            14991: color = 12'h000;
            14992: color = 12'h000;
            14993: color = 12'h000;
            14994: color = 12'h000;
            14995: color = 12'h000;
            14996: color = 12'h000;
            14997: color = 12'h000;
            14998: color = 12'h000;
            14999: color = 12'h000;
            15000: color = 12'h000;
            15001: color = 12'h000;
            15002: color = 12'h000;
            15003: color = 12'h000;
            15004: color = 12'h000;
            15005: color = 12'h000;
            15006: color = 12'h000;
            15007: color = 12'h000;
            15008: color = 12'h000;
            15009: color = 12'h000;
            15010: color = 12'h000;
            15011: color = 12'h000;
            15012: color = 12'h000;
            15013: color = 12'h000;
            15014: color = 12'h000;
            15015: color = 12'h000;
            15016: color = 12'h000;
            15017: color = 12'h000;
            15018: color = 12'h000;
            15019: color = 12'h000;
            15020: color = 12'h000;
            15021: color = 12'h000;
            15022: color = 12'h000;
            15023: color = 12'h000;
            15024: color = 12'h000;
            15025: color = 12'h000;
            15026: color = 12'h000;
            15027: color = 12'h000;
            15028: color = 12'h000;
            15029: color = 12'h000;
            15030: color = 12'h000;
            15031: color = 12'h000;
            15032: color = 12'h000;
            15033: color = 12'h000;
            15034: color = 12'h000;
            15035: color = 12'h000;
            15036: color = 12'h000;
            15037: color = 12'h000;
            15038: color = 12'h000;
            15039: color = 12'h000;
            15040: color = 12'h000;
            15041: color = 12'h000;
            15042: color = 12'h000;
            15043: color = 12'h000;
            15044: color = 12'h000;
            15045: color = 12'h000;
            15046: color = 12'h000;
            15047: color = 12'h000;
            15048: color = 12'h000;
            15049: color = 12'h000;
            15050: color = 12'h000;
            15051: color = 12'h000;
            15052: color = 12'h000;
            15053: color = 12'h000;
            15054: color = 12'h000;
            15055: color = 12'h000;
            15056: color = 12'h000;
            15057: color = 12'h000;
            15058: color = 12'h000;
            15059: color = 12'h000;
            15060: color = 12'h000;
            15061: color = 12'h000;
            15062: color = 12'h000;
            15063: color = 12'h000;
            15064: color = 12'h000;
            15065: color = 12'h000;
            15066: color = 12'h000;
            15067: color = 12'h000;
            15068: color = 12'h000;
            15069: color = 12'h000;
            15070: color = 12'h000;
            15071: color = 12'h000;
            15072: color = 12'h000;
            15073: color = 12'h000;
            15074: color = 12'h000;
            15075: color = 12'h000;
            15076: color = 12'h000;
            15077: color = 12'h000;
            15078: color = 12'h000;
            15079: color = 12'h000;
            15080: color = 12'h000;
            15081: color = 12'h000;
            15082: color = 12'h000;
            15083: color = 12'h000;
            15084: color = 12'h000;
            15085: color = 12'h000;
            15086: color = 12'h000;
            15087: color = 12'h000;
            15088: color = 12'h000;
            15089: color = 12'h000;
            15090: color = 12'h000;
            15091: color = 12'h000;
            15092: color = 12'h000;
            15093: color = 12'h000;
            15094: color = 12'h000;
            15095: color = 12'h000;
            15096: color = 12'h000;
            15097: color = 12'h000;
            15098: color = 12'h000;
            15099: color = 12'h000;
            15100: color = 12'h000;
            15101: color = 12'h000;
            15102: color = 12'h000;
            15103: color = 12'h000;
            15104: color = 12'h000;
            15105: color = 12'h000;
            15106: color = 12'h000;
            15107: color = 12'h000;
            15108: color = 12'h000;
            15109: color = 12'h000;
            15110: color = 12'h000;
            15111: color = 12'h000;
            15112: color = 12'h000;
            15113: color = 12'h000;
            15114: color = 12'h000;
            15115: color = 12'h000;
            15116: color = 12'h000;
            15117: color = 12'h000;
            15118: color = 12'h000;
            15119: color = 12'h000;
            15120: color = 12'h000;
            15121: color = 12'h000;
            15122: color = 12'h000;
            15123: color = 12'h000;
            15124: color = 12'h000;
            15125: color = 12'h000;
            15126: color = 12'h000;
            15127: color = 12'h000;
            15128: color = 12'h000;
            15129: color = 12'h000;
            15130: color = 12'h000;
            15131: color = 12'h000;
            15132: color = 12'h000;
            15133: color = 12'h000;
            15134: color = 12'h000;
            15135: color = 12'h000;
            15136: color = 12'h000;
            15137: color = 12'h000;
            15138: color = 12'h000;
            15139: color = 12'h000;
            15140: color = 12'h000;
            15141: color = 12'h000;
            15142: color = 12'h000;
            15143: color = 12'h000;
            15144: color = 12'h000;
            15145: color = 12'h000;
            15146: color = 12'h000;
            15147: color = 12'h000;
            15148: color = 12'h000;
            15149: color = 12'h000;
            15150: color = 12'h000;
            15151: color = 12'h000;
            15152: color = 12'h000;
            15153: color = 12'h000;
            15154: color = 12'h000;
            15155: color = 12'h000;
            15156: color = 12'h000;
            15157: color = 12'h000;
            15158: color = 12'h000;
            15159: color = 12'h000;
            15160: color = 12'h000;
            15161: color = 12'h000;
            15162: color = 12'h000;
            15163: color = 12'h000;
            15164: color = 12'h000;
            15165: color = 12'h000;
            15166: color = 12'h000;
            15167: color = 12'h000;
            15168: color = 12'h000;
            15169: color = 12'h000;
            15170: color = 12'h000;
            15171: color = 12'h000;
            15172: color = 12'h000;
            15173: color = 12'h000;
            15174: color = 12'h000;
            15175: color = 12'h000;
            15176: color = 12'h000;
            15177: color = 12'h000;
            15178: color = 12'h000;
            15179: color = 12'h000;
            15180: color = 12'h000;
            15181: color = 12'h000;
            15182: color = 12'h000;
            15183: color = 12'h000;
            15184: color = 12'h000;
            15185: color = 12'h000;
            15186: color = 12'h000;
            15187: color = 12'h000;
            15188: color = 12'h000;
            15189: color = 12'h000;
            15190: color = 12'h000;
            15191: color = 12'h000;
            15192: color = 12'h000;
            15193: color = 12'h000;
            15194: color = 12'h000;
            15195: color = 12'h000;
            15196: color = 12'h000;
            15197: color = 12'h000;
            15198: color = 12'h000;
            15199: color = 12'h000;
            15200: color = 12'h000;
            15201: color = 12'h000;
            15202: color = 12'h000;
            15203: color = 12'h000;
            15204: color = 12'h000;
            15205: color = 12'h000;
            15206: color = 12'h000;
            15207: color = 12'h000;
            15208: color = 12'h000;
            15209: color = 12'h000;
            15210: color = 12'h000;
            15211: color = 12'h000;
            15212: color = 12'h000;
            15213: color = 12'h000;
            15214: color = 12'h000;
            15215: color = 12'h000;
            15216: color = 12'h000;
            15217: color = 12'h000;
            15218: color = 12'h000;
            15219: color = 12'h000;
            15220: color = 12'h000;
            15221: color = 12'h000;
            15222: color = 12'h000;
            15223: color = 12'h000;
            15224: color = 12'h000;
            15225: color = 12'h000;
            15226: color = 12'h000;
            15227: color = 12'h000;
            15228: color = 12'h000;
            15229: color = 12'h000;
            15230: color = 12'h000;
            15231: color = 12'h000;
            15232: color = 12'h000;
            15233: color = 12'h000;
            15234: color = 12'h000;
            15235: color = 12'h000;
            15236: color = 12'h000;
            15237: color = 12'h000;
            15238: color = 12'h000;
            15239: color = 12'h000;
            15240: color = 12'h000;
            15241: color = 12'h000;
            15242: color = 12'h000;
            15243: color = 12'h000;
            15244: color = 12'h000;
            15245: color = 12'h000;
            15246: color = 12'h000;
            15247: color = 12'h000;
            15248: color = 12'h000;
            15249: color = 12'h000;
            15250: color = 12'h000;
            15251: color = 12'h000;
            15252: color = 12'h000;
            15253: color = 12'h000;
            15254: color = 12'h000;
            15255: color = 12'h000;
            15256: color = 12'h000;
            15257: color = 12'h000;
            15258: color = 12'h000;
            15259: color = 12'h000;
            15260: color = 12'h000;
            15261: color = 12'h000;
            15262: color = 12'h000;
            15263: color = 12'h000;
            15264: color = 12'h000;
            15265: color = 12'h000;
            15266: color = 12'h000;
            15267: color = 12'h000;
            15268: color = 12'h000;
            15269: color = 12'h000;
            15270: color = 12'h000;
            15271: color = 12'h000;
            15272: color = 12'h000;
            15273: color = 12'h000;
            15274: color = 12'h000;
            15275: color = 12'h000;
            15276: color = 12'h000;
            15277: color = 12'h000;
            15278: color = 12'h000;
            15279: color = 12'h000;
            15280: color = 12'h000;
            15281: color = 12'h000;
            15282: color = 12'h000;
            15283: color = 12'h000;
            15284: color = 12'h000;
            15285: color = 12'h000;
            15286: color = 12'h000;
            15287: color = 12'h000;
            15288: color = 12'h000;
            15289: color = 12'h000;
            15290: color = 12'h000;
            15291: color = 12'h000;
            15292: color = 12'h000;
            15293: color = 12'h000;
            15294: color = 12'h000;
            15295: color = 12'h000;
            15296: color = 12'h000;
            15297: color = 12'h000;
            15298: color = 12'h000;
            15299: color = 12'h000;
            15300: color = 12'h000;
            15301: color = 12'h000;
            15302: color = 12'h000;
            15303: color = 12'h000;
            15304: color = 12'h000;
            15305: color = 12'h000;
            15306: color = 12'h000;
            15307: color = 12'h000;
            15308: color = 12'h000;
            15309: color = 12'h000;
            15310: color = 12'h000;
            15311: color = 12'h000;
            15312: color = 12'h000;
            15313: color = 12'h000;
            15314: color = 12'h000;
            15315: color = 12'h000;
            15316: color = 12'h000;
            15317: color = 12'h000;
            15318: color = 12'h000;
            15319: color = 12'h000;
            15320: color = 12'h000;
            15321: color = 12'h000;
            15322: color = 12'h000;
            15323: color = 12'h000;
            15324: color = 12'h000;
            15325: color = 12'h000;
            15326: color = 12'h000;
            15327: color = 12'h000;
            15328: color = 12'h000;
            15329: color = 12'h000;
            15330: color = 12'h000;
            15331: color = 12'h000;
            15332: color = 12'h000;
            15333: color = 12'h000;
            15334: color = 12'h000;
            15335: color = 12'h000;
            15336: color = 12'h000;
            15337: color = 12'h000;
            15338: color = 12'h000;
            15339: color = 12'h000;
            15340: color = 12'h000;
            15341: color = 12'h000;
            15342: color = 12'h000;
            15343: color = 12'h000;
            15344: color = 12'h000;
            15345: color = 12'h000;
            15346: color = 12'h000;
            15347: color = 12'h000;
            15348: color = 12'h000;
            15349: color = 12'h000;
            15350: color = 12'h000;
            15351: color = 12'h000;
            15352: color = 12'h000;
            15353: color = 12'h000;
            15354: color = 12'h000;
            15355: color = 12'h000;
            15356: color = 12'h000;
            15357: color = 12'h000;
            15358: color = 12'h000;
            15359: color = 12'h000;
            15360: color = 12'h000;
            15361: color = 12'h000;
            15362: color = 12'h000;
            15363: color = 12'h000;
            15364: color = 12'h000;
            15365: color = 12'h000;
            15366: color = 12'h000;
            15367: color = 12'h000;
            15368: color = 12'h000;
            15369: color = 12'h000;
            15370: color = 12'h000;
            15371: color = 12'h000;
            15372: color = 12'h000;
            15373: color = 12'h000;
            15374: color = 12'h000;
            15375: color = 12'h000;
            15376: color = 12'h000;
            15377: color = 12'h000;
            15378: color = 12'h000;
            15379: color = 12'h000;
            15380: color = 12'h000;
            15381: color = 12'h000;
            15382: color = 12'h000;
            15383: color = 12'h000;
            15384: color = 12'h000;
            15385: color = 12'h000;
            15386: color = 12'h000;
            15387: color = 12'h000;
            15388: color = 12'h000;
            15389: color = 12'h000;
            15390: color = 12'h000;
            15391: color = 12'h000;
            15392: color = 12'h000;
            15393: color = 12'h000;
            15394: color = 12'h000;
            15395: color = 12'h000;
            15396: color = 12'h000;
            15397: color = 12'h000;
            15398: color = 12'h000;
            15399: color = 12'h000;
            15400: color = 12'h000;
            15401: color = 12'h000;
            15402: color = 12'h000;
            15403: color = 12'h000;
            15404: color = 12'h000;
            15405: color = 12'h000;
            15406: color = 12'h000;
            15407: color = 12'h000;
            15408: color = 12'h000;
            15409: color = 12'h000;
            15410: color = 12'h000;
            15411: color = 12'h000;
            15412: color = 12'h000;
            15413: color = 12'h000;
            15414: color = 12'h000;
            15415: color = 12'h000;
            15416: color = 12'h000;
            15417: color = 12'h000;
            15418: color = 12'h000;
            15419: color = 12'h000;
            15420: color = 12'h000;
            15421: color = 12'h000;
            15422: color = 12'h000;
            15423: color = 12'h000;
            15424: color = 12'h000;
            15425: color = 12'h000;
            15426: color = 12'h000;
            15427: color = 12'h000;
            15428: color = 12'h000;
            15429: color = 12'h000;
            15430: color = 12'h000;
            15431: color = 12'h000;
            15432: color = 12'h000;
            15433: color = 12'h000;
            15434: color = 12'h000;
            15435: color = 12'h000;
            15436: color = 12'h000;
            15437: color = 12'h000;
            15438: color = 12'h000;
            15439: color = 12'h000;
            15440: color = 12'h000;
            15441: color = 12'h000;
            15442: color = 12'h000;
            15443: color = 12'h000;
            15444: color = 12'h000;
            15445: color = 12'h000;
            15446: color = 12'h000;
            15447: color = 12'h000;
            15448: color = 12'h000;
            15449: color = 12'h000;
            15450: color = 12'h000;
            15451: color = 12'h000;
            15452: color = 12'h000;
            15453: color = 12'h000;
            15454: color = 12'h000;
            15455: color = 12'h000;
            15456: color = 12'h000;
            15457: color = 12'h000;
            15458: color = 12'h000;
            15459: color = 12'h000;
            15460: color = 12'h000;
            15461: color = 12'h000;
            15462: color = 12'h000;
            15463: color = 12'h000;
            15464: color = 12'h000;
            15465: color = 12'h000;
            15466: color = 12'h000;
            15467: color = 12'h000;
            15468: color = 12'h000;
            15469: color = 12'h000;
            15470: color = 12'h000;
            15471: color = 12'h000;
            15472: color = 12'h000;
            15473: color = 12'h000;
            15474: color = 12'h000;
            15475: color = 12'h000;
            15476: color = 12'h000;
            15477: color = 12'h000;
            15478: color = 12'h000;
            15479: color = 12'h000;
            15480: color = 12'h000;
            15481: color = 12'h000;
            15482: color = 12'h000;
            15483: color = 12'h000;
            15484: color = 12'h000;
            15485: color = 12'h000;
            15486: color = 12'h000;
            15487: color = 12'h000;
            15488: color = 12'h000;
            15489: color = 12'h000;
            15490: color = 12'h000;
            15491: color = 12'h000;
            15492: color = 12'h000;
            15493: color = 12'h000;
            15494: color = 12'h000;
            15495: color = 12'h000;
            15496: color = 12'h000;
            15497: color = 12'h000;
            15498: color = 12'h000;
            15499: color = 12'h000;
            15500: color = 12'h000;
            15501: color = 12'h000;
            15502: color = 12'h000;
            15503: color = 12'h000;
            15504: color = 12'h000;
            15505: color = 12'h000;
            15506: color = 12'h000;
            15507: color = 12'h000;
            15508: color = 12'h000;
            15509: color = 12'h000;
            15510: color = 12'h000;
            15511: color = 12'h000;
            15512: color = 12'h000;
            15513: color = 12'h000;
            15514: color = 12'h000;
            15515: color = 12'h000;
            15516: color = 12'h000;
            15517: color = 12'h000;
            15518: color = 12'h000;
            15519: color = 12'h000;
            15520: color = 12'h000;
            15521: color = 12'h000;
            15522: color = 12'h000;
            15523: color = 12'h000;
            15524: color = 12'h000;
            15525: color = 12'h000;
            15526: color = 12'h000;
            15527: color = 12'h000;
            15528: color = 12'h000;
            15529: color = 12'h000;
            15530: color = 12'h000;
            15531: color = 12'h000;
            15532: color = 12'h000;
            15533: color = 12'h000;
            15534: color = 12'h000;
            15535: color = 12'h000;
            15536: color = 12'h000;
            15537: color = 12'h000;
            15538: color = 12'h000;
            15539: color = 12'h000;
            15540: color = 12'h000;
            15541: color = 12'h000;
            15542: color = 12'h000;
            15543: color = 12'h000;
            15544: color = 12'h000;
            15545: color = 12'h000;
            15546: color = 12'h000;
            15547: color = 12'h000;
            15548: color = 12'h000;
            15549: color = 12'h000;
            15550: color = 12'h000;
            15551: color = 12'h000;
            15552: color = 12'h000;
            15553: color = 12'h000;
            15554: color = 12'h000;
            15555: color = 12'h000;
            15556: color = 12'h000;
            15557: color = 12'h000;
            15558: color = 12'h000;
            15559: color = 12'h000;
            15560: color = 12'h000;
            15561: color = 12'h000;
            15562: color = 12'h000;
            15563: color = 12'h000;
            15564: color = 12'h000;
            15565: color = 12'h000;
            15566: color = 12'h000;
            15567: color = 12'h000;
            15568: color = 12'h000;
            15569: color = 12'h000;
            15570: color = 12'h000;
            15571: color = 12'h000;
            15572: color = 12'h000;
            15573: color = 12'h000;
            15574: color = 12'h000;
            15575: color = 12'h000;
            15576: color = 12'h000;
            15577: color = 12'h000;
            15578: color = 12'h000;
            15579: color = 12'h000;
            15580: color = 12'h000;
            15581: color = 12'h000;
            15582: color = 12'h000;
            15583: color = 12'h000;
            15584: color = 12'h000;
            15585: color = 12'h000;
            15586: color = 12'h000;
            15587: color = 12'h000;
            15588: color = 12'h000;
            15589: color = 12'h000;
            15590: color = 12'h000;
            15591: color = 12'h000;
            15592: color = 12'h000;
            15593: color = 12'h000;
            15594: color = 12'h000;
            15595: color = 12'h000;
            15596: color = 12'h000;
            15597: color = 12'h000;
            15598: color = 12'h000;
            15599: color = 12'h000;
            15600: color = 12'h000;
            15601: color = 12'h000;
            15602: color = 12'h000;
            15603: color = 12'h000;
            15604: color = 12'h000;
            15605: color = 12'h000;
            15606: color = 12'h000;
            15607: color = 12'h000;
            15608: color = 12'h000;
            15609: color = 12'h000;
            15610: color = 12'h000;
            15611: color = 12'h000;
            15612: color = 12'h000;
            15613: color = 12'h000;
            15614: color = 12'h000;
            15615: color = 12'h000;
            15616: color = 12'h000;
            15617: color = 12'h000;
            15618: color = 12'h000;
            15619: color = 12'h000;
            15620: color = 12'h000;
            15621: color = 12'h000;
            15622: color = 12'h000;
            15623: color = 12'h000;
            15624: color = 12'h000;
            15625: color = 12'h000;
            15626: color = 12'h000;
            15627: color = 12'h000;
            15628: color = 12'h000;
            15629: color = 12'h000;
            15630: color = 12'h000;
            15631: color = 12'h000;
            15632: color = 12'h000;
            15633: color = 12'h000;
            15634: color = 12'h000;
            15635: color = 12'h000;
            15636: color = 12'h000;
            15637: color = 12'h000;
            15638: color = 12'h000;
            15639: color = 12'h000;
            15640: color = 12'h000;
            15641: color = 12'h000;
            15642: color = 12'h000;
            15643: color = 12'h000;
            15644: color = 12'h000;
            15645: color = 12'h000;
            15646: color = 12'h000;
            15647: color = 12'h000;
            15648: color = 12'h000;
            15649: color = 12'h000;
            15650: color = 12'h000;
            15651: color = 12'h000;
            15652: color = 12'h000;
            15653: color = 12'h000;
            15654: color = 12'h000;
            15655: color = 12'h000;
            15656: color = 12'h000;
            15657: color = 12'h000;
            15658: color = 12'h000;
            15659: color = 12'h000;
            15660: color = 12'h000;
            15661: color = 12'h000;
            15662: color = 12'h000;
            15663: color = 12'h000;
            15664: color = 12'h000;
            15665: color = 12'h000;
            15666: color = 12'h000;
            15667: color = 12'h000;
            15668: color = 12'h000;
            15669: color = 12'h000;
            15670: color = 12'h000;
            15671: color = 12'h000;
            15672: color = 12'h000;
            15673: color = 12'h000;
            15674: color = 12'h000;
            15675: color = 12'h000;
            15676: color = 12'h000;
            15677: color = 12'h000;
            15678: color = 12'h000;
            15679: color = 12'h000;
            15680: color = 12'h000;
            15681: color = 12'h000;
            15682: color = 12'h000;
            15683: color = 12'h000;
            15684: color = 12'h000;
            15685: color = 12'h000;
            15686: color = 12'h000;
            15687: color = 12'h000;
            15688: color = 12'h000;
            15689: color = 12'h000;
            15690: color = 12'h000;
            15691: color = 12'h000;
            15692: color = 12'h000;
            15693: color = 12'h000;
            15694: color = 12'h000;
            15695: color = 12'h000;
            15696: color = 12'h000;
            15697: color = 12'h000;
            15698: color = 12'h000;
            15699: color = 12'h000;
            15700: color = 12'h000;
            15701: color = 12'h000;
            15702: color = 12'h000;
            15703: color = 12'h000;
            15704: color = 12'h000;
            15705: color = 12'h000;
            15706: color = 12'h000;
            15707: color = 12'h000;
            15708: color = 12'h000;
            15709: color = 12'h000;
            15710: color = 12'h000;
            15711: color = 12'h000;
            15712: color = 12'h000;
            15713: color = 12'h000;
            15714: color = 12'h000;
            15715: color = 12'h000;
            15716: color = 12'h000;
            15717: color = 12'h000;
            15718: color = 12'h000;
            15719: color = 12'h000;
            15720: color = 12'h000;
            15721: color = 12'h000;
            15722: color = 12'h000;
            15723: color = 12'h000;
            15724: color = 12'h000;
            15725: color = 12'h000;
            15726: color = 12'h000;
            15727: color = 12'h000;
            15728: color = 12'h000;
            15729: color = 12'h000;
            15730: color = 12'h000;
            15731: color = 12'h000;
            15732: color = 12'h000;
            15733: color = 12'h000;
            15734: color = 12'h000;
            15735: color = 12'h000;
            15736: color = 12'h000;
            15737: color = 12'h000;
            15738: color = 12'h000;
            15739: color = 12'h000;
            15740: color = 12'h000;
            15741: color = 12'h000;
            15742: color = 12'h000;
            15743: color = 12'h000;
            15744: color = 12'h000;
            15745: color = 12'h000;
            15746: color = 12'h000;
            15747: color = 12'h000;
            15748: color = 12'h000;
            15749: color = 12'h000;
            15750: color = 12'h000;
            15751: color = 12'h000;
            15752: color = 12'h000;
            15753: color = 12'h000;
            15754: color = 12'h000;
            15755: color = 12'h000;
            15756: color = 12'h000;
            15757: color = 12'h000;
            15758: color = 12'h000;
            15759: color = 12'h000;
            15760: color = 12'h000;
            15761: color = 12'h000;
            15762: color = 12'h000;
            15763: color = 12'h000;
            15764: color = 12'h000;
            15765: color = 12'h000;
            15766: color = 12'h000;
            15767: color = 12'h000;
            15768: color = 12'h000;
            15769: color = 12'h000;
            15770: color = 12'h000;
            15771: color = 12'h000;
            15772: color = 12'h000;
            15773: color = 12'h000;
            15774: color = 12'h000;
            15775: color = 12'h000;
            15776: color = 12'h000;
            15777: color = 12'h000;
            15778: color = 12'h000;
            15779: color = 12'h000;
            15780: color = 12'h000;
            15781: color = 12'h000;
            15782: color = 12'h000;
            15783: color = 12'h000;
            15784: color = 12'h000;
            15785: color = 12'h000;
            15786: color = 12'h000;
            15787: color = 12'h000;
            15788: color = 12'h000;
            15789: color = 12'h000;
            15790: color = 12'h000;
            15791: color = 12'h000;
            15792: color = 12'h000;
            15793: color = 12'h000;
            15794: color = 12'h000;
            15795: color = 12'h000;
            15796: color = 12'h000;
            15797: color = 12'h000;
            15798: color = 12'h000;
            15799: color = 12'h000;
            15800: color = 12'h000;
            15801: color = 12'h000;
            15802: color = 12'h000;
            15803: color = 12'h000;
            15804: color = 12'h000;
            15805: color = 12'h000;
            15806: color = 12'h000;
            15807: color = 12'h000;
            15808: color = 12'h000;
            15809: color = 12'h000;
            15810: color = 12'h000;
            15811: color = 12'h000;
            15812: color = 12'h000;
            15813: color = 12'h000;
            15814: color = 12'h000;
            15815: color = 12'h000;
            15816: color = 12'h000;
            15817: color = 12'h000;
            15818: color = 12'h000;
            15819: color = 12'h000;
            15820: color = 12'h000;
            15821: color = 12'h000;
            15822: color = 12'h000;
            15823: color = 12'h000;
            15824: color = 12'h000;
            15825: color = 12'h000;
            15826: color = 12'h000;
            15827: color = 12'h000;
            15828: color = 12'h000;
            15829: color = 12'h000;
            15830: color = 12'h000;
            15831: color = 12'h000;
            15832: color = 12'h000;
            15833: color = 12'h000;
            15834: color = 12'h000;
            15835: color = 12'h000;
            15836: color = 12'h000;
            15837: color = 12'h000;
            15838: color = 12'h000;
            15839: color = 12'h000;
            15840: color = 12'h000;
            15841: color = 12'h000;
            15842: color = 12'h000;
            15843: color = 12'h000;
            15844: color = 12'h000;
            15845: color = 12'h000;
            15846: color = 12'h000;
            15847: color = 12'h000;
            15848: color = 12'h000;
            15849: color = 12'h000;
            15850: color = 12'h000;
            15851: color = 12'h000;
            15852: color = 12'h000;
            15853: color = 12'h000;
            15854: color = 12'h000;
            15855: color = 12'h000;
            15856: color = 12'h000;
            15857: color = 12'h000;
            15858: color = 12'h000;
            15859: color = 12'h000;
            15860: color = 12'h000;
            15861: color = 12'h000;
            15862: color = 12'h000;
            15863: color = 12'h000;
            15864: color = 12'h000;
            15865: color = 12'h000;
            15866: color = 12'h000;
            15867: color = 12'h000;
            15868: color = 12'h000;
            15869: color = 12'h000;
            15870: color = 12'h000;
            15871: color = 12'h000;
            15872: color = 12'h000;
            15873: color = 12'h000;
            15874: color = 12'h000;
            15875: color = 12'h000;
            15876: color = 12'h000;
            15877: color = 12'h000;
            15878: color = 12'h000;
            15879: color = 12'h000;
            15880: color = 12'h000;
            15881: color = 12'h000;
            15882: color = 12'h000;
            15883: color = 12'h000;
            15884: color = 12'h000;
            15885: color = 12'h000;
            15886: color = 12'h000;
            15887: color = 12'h000;
            15888: color = 12'h000;
            15889: color = 12'h000;
            15890: color = 12'h000;
            15891: color = 12'h000;
            15892: color = 12'h000;
            15893: color = 12'h000;
            15894: color = 12'h000;
            15895: color = 12'h000;
            15896: color = 12'h000;
            15897: color = 12'h000;
            15898: color = 12'h000;
            15899: color = 12'h000;
            15900: color = 12'h000;
            15901: color = 12'h000;
            15902: color = 12'h000;
            15903: color = 12'h000;
            15904: color = 12'h000;
            15905: color = 12'h000;
            15906: color = 12'h000;
            15907: color = 12'h000;
            15908: color = 12'h000;
            15909: color = 12'h000;
            15910: color = 12'h000;
            15911: color = 12'h000;
            15912: color = 12'h000;
            15913: color = 12'h000;
            15914: color = 12'h000;
            15915: color = 12'h000;
            15916: color = 12'h000;
            15917: color = 12'h000;
            15918: color = 12'h000;
            15919: color = 12'h000;
            15920: color = 12'h000;
            15921: color = 12'h000;
            15922: color = 12'h000;
            15923: color = 12'h000;
            15924: color = 12'h000;
            15925: color = 12'h000;
            15926: color = 12'h000;
            15927: color = 12'h000;
            15928: color = 12'h000;
            15929: color = 12'h000;
            15930: color = 12'h000;
            15931: color = 12'h000;
            15932: color = 12'h000;
            15933: color = 12'h000;
            15934: color = 12'h000;
            15935: color = 12'h000;
            15936: color = 12'h000;
            15937: color = 12'h000;
            15938: color = 12'h000;
            15939: color = 12'h000;
            15940: color = 12'h000;
            15941: color = 12'h000;
            15942: color = 12'h000;
            15943: color = 12'h000;
            15944: color = 12'h000;
            15945: color = 12'h000;
            15946: color = 12'h000;
            15947: color = 12'h000;
            15948: color = 12'h000;
            15949: color = 12'h000;
            15950: color = 12'h000;
            15951: color = 12'h000;
            15952: color = 12'h000;
            15953: color = 12'h000;
            15954: color = 12'h000;
            15955: color = 12'h000;
            15956: color = 12'h000;
            15957: color = 12'h000;
            15958: color = 12'h000;
            15959: color = 12'h000;
            15960: color = 12'h000;
            15961: color = 12'h000;
            15962: color = 12'h000;
            15963: color = 12'h000;
            15964: color = 12'h000;
            15965: color = 12'h000;
            15966: color = 12'h000;
            15967: color = 12'h000;
            15968: color = 12'h000;
            15969: color = 12'h000;
            15970: color = 12'h000;
            15971: color = 12'h000;
            15972: color = 12'h000;
            15973: color = 12'h000;
            15974: color = 12'h000;
            15975: color = 12'h000;
            15976: color = 12'h000;
            15977: color = 12'h000;
            15978: color = 12'h000;
            15979: color = 12'h000;
            15980: color = 12'h000;
            15981: color = 12'h000;
            15982: color = 12'h000;
            15983: color = 12'h000;
            15984: color = 12'h000;
            15985: color = 12'h000;
            15986: color = 12'h000;
            15987: color = 12'h000;
            15988: color = 12'h000;
            15989: color = 12'h000;
            15990: color = 12'h000;
            15991: color = 12'h000;
            15992: color = 12'h000;
            15993: color = 12'h000;
            15994: color = 12'h000;
            15995: color = 12'h000;
            15996: color = 12'h000;
            15997: color = 12'h000;
            15998: color = 12'h000;
            15999: color = 12'h000;
            default: color = 12'h000;
        endcase
    end
endmodule